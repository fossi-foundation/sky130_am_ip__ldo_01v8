magic
tech sky130A
timestamp 1713186496
<< pwell >>
rect -139 -10129 139 10129
<< mvnmos >>
rect -25 -10000 25 10000
<< mvndiff >>
rect -54 9994 -25 10000
rect -54 -9994 -48 9994
rect -31 -9994 -25 9994
rect -54 -10000 -25 -9994
rect 25 9994 54 10000
rect 25 -9994 31 9994
rect 48 -9994 54 9994
rect 25 -10000 54 -9994
<< mvndiffc >>
rect -48 -9994 -31 9994
rect 31 -9994 48 9994
<< mvpsubdiff >>
rect -121 10105 121 10111
rect -121 10088 -67 10105
rect 67 10088 121 10105
rect -121 10082 121 10088
rect -121 10057 -92 10082
rect -121 -10057 -115 10057
rect -98 -10057 -92 10057
rect 92 10057 121 10082
rect -121 -10082 -92 -10057
rect 92 -10057 98 10057
rect 115 -10057 121 10057
rect 92 -10082 121 -10057
rect -121 -10088 121 -10082
rect -121 -10105 -67 -10088
rect 67 -10105 121 -10088
rect -121 -10111 121 -10105
<< mvpsubdiffcont >>
rect -67 10088 67 10105
rect -115 -10057 -98 10057
rect 98 -10057 115 10057
rect -67 -10105 67 -10088
<< poly >>
rect -25 10036 25 10044
rect -25 10019 -17 10036
rect 17 10019 25 10036
rect -25 10000 25 10019
rect -25 -10019 25 -10000
rect -25 -10036 -17 -10019
rect 17 -10036 25 -10019
rect -25 -10044 25 -10036
<< polycont >>
rect -17 10019 17 10036
rect -17 -10036 17 -10019
<< locali >>
rect -115 10088 -67 10105
rect 67 10088 115 10105
rect -115 10057 -98 10088
rect 98 10057 115 10088
rect -25 10019 -17 10036
rect 17 10019 25 10036
rect -48 9994 -31 10002
rect -48 -10002 -31 -9994
rect 31 9994 48 10002
rect 31 -10002 48 -9994
rect -25 -10036 -17 -10019
rect 17 -10036 25 -10019
rect -115 -10088 -98 -10057
rect 98 -10088 115 -10057
rect -115 -10105 -67 -10088
rect 67 -10105 115 -10088
<< viali >>
rect -17 10019 17 10036
rect -48 -9994 -31 9994
rect 31 -9994 48 9994
rect -17 -10036 17 -10019
<< metal1 >>
rect -23 10036 23 10039
rect -23 10019 -17 10036
rect 17 10019 23 10036
rect -23 10016 23 10019
rect -51 9994 -28 10000
rect -51 -9994 -48 9994
rect -31 -9994 -28 9994
rect -51 -10000 -28 -9994
rect 28 9994 51 10000
rect 28 -9994 31 9994
rect 48 -9994 51 9994
rect 28 -10000 51 -9994
rect -23 -10019 23 -10016
rect -23 -10036 -17 -10019
rect 17 -10036 23 -10019
rect -23 -10039 23 -10036
<< properties >>
string FIXED_BBOX -106 -10096 106 10096
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 200.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
