magic
tech sky130A
magscale 1 2
timestamp 1726591810
<< pwell >>
rect -1789 -6239 1789 6239
<< mvnmos >>
rect -1551 4981 -1451 5981
rect -1393 4981 -1293 5981
rect -1235 4981 -1135 5981
rect -1077 4981 -977 5981
rect -919 4981 -819 5981
rect -761 4981 -661 5981
rect -603 4981 -503 5981
rect -445 4981 -345 5981
rect -287 4981 -187 5981
rect -129 4981 -29 5981
rect 29 4981 129 5981
rect 187 4981 287 5981
rect 345 4981 445 5981
rect 503 4981 603 5981
rect 661 4981 761 5981
rect 819 4981 919 5981
rect 977 4981 1077 5981
rect 1135 4981 1235 5981
rect 1293 4981 1393 5981
rect 1451 4981 1551 5981
rect -1551 3763 -1451 4763
rect -1393 3763 -1293 4763
rect -1235 3763 -1135 4763
rect -1077 3763 -977 4763
rect -919 3763 -819 4763
rect -761 3763 -661 4763
rect -603 3763 -503 4763
rect -445 3763 -345 4763
rect -287 3763 -187 4763
rect -129 3763 -29 4763
rect 29 3763 129 4763
rect 187 3763 287 4763
rect 345 3763 445 4763
rect 503 3763 603 4763
rect 661 3763 761 4763
rect 819 3763 919 4763
rect 977 3763 1077 4763
rect 1135 3763 1235 4763
rect 1293 3763 1393 4763
rect 1451 3763 1551 4763
rect -1551 2545 -1451 3545
rect -1393 2545 -1293 3545
rect -1235 2545 -1135 3545
rect -1077 2545 -977 3545
rect -919 2545 -819 3545
rect -761 2545 -661 3545
rect -603 2545 -503 3545
rect -445 2545 -345 3545
rect -287 2545 -187 3545
rect -129 2545 -29 3545
rect 29 2545 129 3545
rect 187 2545 287 3545
rect 345 2545 445 3545
rect 503 2545 603 3545
rect 661 2545 761 3545
rect 819 2545 919 3545
rect 977 2545 1077 3545
rect 1135 2545 1235 3545
rect 1293 2545 1393 3545
rect 1451 2545 1551 3545
rect -1551 1327 -1451 2327
rect -1393 1327 -1293 2327
rect -1235 1327 -1135 2327
rect -1077 1327 -977 2327
rect -919 1327 -819 2327
rect -761 1327 -661 2327
rect -603 1327 -503 2327
rect -445 1327 -345 2327
rect -287 1327 -187 2327
rect -129 1327 -29 2327
rect 29 1327 129 2327
rect 187 1327 287 2327
rect 345 1327 445 2327
rect 503 1327 603 2327
rect 661 1327 761 2327
rect 819 1327 919 2327
rect 977 1327 1077 2327
rect 1135 1327 1235 2327
rect 1293 1327 1393 2327
rect 1451 1327 1551 2327
rect -1551 109 -1451 1109
rect -1393 109 -1293 1109
rect -1235 109 -1135 1109
rect -1077 109 -977 1109
rect -919 109 -819 1109
rect -761 109 -661 1109
rect -603 109 -503 1109
rect -445 109 -345 1109
rect -287 109 -187 1109
rect -129 109 -29 1109
rect 29 109 129 1109
rect 187 109 287 1109
rect 345 109 445 1109
rect 503 109 603 1109
rect 661 109 761 1109
rect 819 109 919 1109
rect 977 109 1077 1109
rect 1135 109 1235 1109
rect 1293 109 1393 1109
rect 1451 109 1551 1109
rect -1551 -1109 -1451 -109
rect -1393 -1109 -1293 -109
rect -1235 -1109 -1135 -109
rect -1077 -1109 -977 -109
rect -919 -1109 -819 -109
rect -761 -1109 -661 -109
rect -603 -1109 -503 -109
rect -445 -1109 -345 -109
rect -287 -1109 -187 -109
rect -129 -1109 -29 -109
rect 29 -1109 129 -109
rect 187 -1109 287 -109
rect 345 -1109 445 -109
rect 503 -1109 603 -109
rect 661 -1109 761 -109
rect 819 -1109 919 -109
rect 977 -1109 1077 -109
rect 1135 -1109 1235 -109
rect 1293 -1109 1393 -109
rect 1451 -1109 1551 -109
rect -1551 -2327 -1451 -1327
rect -1393 -2327 -1293 -1327
rect -1235 -2327 -1135 -1327
rect -1077 -2327 -977 -1327
rect -919 -2327 -819 -1327
rect -761 -2327 -661 -1327
rect -603 -2327 -503 -1327
rect -445 -2327 -345 -1327
rect -287 -2327 -187 -1327
rect -129 -2327 -29 -1327
rect 29 -2327 129 -1327
rect 187 -2327 287 -1327
rect 345 -2327 445 -1327
rect 503 -2327 603 -1327
rect 661 -2327 761 -1327
rect 819 -2327 919 -1327
rect 977 -2327 1077 -1327
rect 1135 -2327 1235 -1327
rect 1293 -2327 1393 -1327
rect 1451 -2327 1551 -1327
rect -1551 -3545 -1451 -2545
rect -1393 -3545 -1293 -2545
rect -1235 -3545 -1135 -2545
rect -1077 -3545 -977 -2545
rect -919 -3545 -819 -2545
rect -761 -3545 -661 -2545
rect -603 -3545 -503 -2545
rect -445 -3545 -345 -2545
rect -287 -3545 -187 -2545
rect -129 -3545 -29 -2545
rect 29 -3545 129 -2545
rect 187 -3545 287 -2545
rect 345 -3545 445 -2545
rect 503 -3545 603 -2545
rect 661 -3545 761 -2545
rect 819 -3545 919 -2545
rect 977 -3545 1077 -2545
rect 1135 -3545 1235 -2545
rect 1293 -3545 1393 -2545
rect 1451 -3545 1551 -2545
rect -1551 -4763 -1451 -3763
rect -1393 -4763 -1293 -3763
rect -1235 -4763 -1135 -3763
rect -1077 -4763 -977 -3763
rect -919 -4763 -819 -3763
rect -761 -4763 -661 -3763
rect -603 -4763 -503 -3763
rect -445 -4763 -345 -3763
rect -287 -4763 -187 -3763
rect -129 -4763 -29 -3763
rect 29 -4763 129 -3763
rect 187 -4763 287 -3763
rect 345 -4763 445 -3763
rect 503 -4763 603 -3763
rect 661 -4763 761 -3763
rect 819 -4763 919 -3763
rect 977 -4763 1077 -3763
rect 1135 -4763 1235 -3763
rect 1293 -4763 1393 -3763
rect 1451 -4763 1551 -3763
rect -1551 -5981 -1451 -4981
rect -1393 -5981 -1293 -4981
rect -1235 -5981 -1135 -4981
rect -1077 -5981 -977 -4981
rect -919 -5981 -819 -4981
rect -761 -5981 -661 -4981
rect -603 -5981 -503 -4981
rect -445 -5981 -345 -4981
rect -287 -5981 -187 -4981
rect -129 -5981 -29 -4981
rect 29 -5981 129 -4981
rect 187 -5981 287 -4981
rect 345 -5981 445 -4981
rect 503 -5981 603 -4981
rect 661 -5981 761 -4981
rect 819 -5981 919 -4981
rect 977 -5981 1077 -4981
rect 1135 -5981 1235 -4981
rect 1293 -5981 1393 -4981
rect 1451 -5981 1551 -4981
<< mvndiff >>
rect -1609 5969 -1551 5981
rect -1609 4993 -1597 5969
rect -1563 4993 -1551 5969
rect -1609 4981 -1551 4993
rect -1451 5969 -1393 5981
rect -1451 4993 -1439 5969
rect -1405 4993 -1393 5969
rect -1451 4981 -1393 4993
rect -1293 5969 -1235 5981
rect -1293 4993 -1281 5969
rect -1247 4993 -1235 5969
rect -1293 4981 -1235 4993
rect -1135 5969 -1077 5981
rect -1135 4993 -1123 5969
rect -1089 4993 -1077 5969
rect -1135 4981 -1077 4993
rect -977 5969 -919 5981
rect -977 4993 -965 5969
rect -931 4993 -919 5969
rect -977 4981 -919 4993
rect -819 5969 -761 5981
rect -819 4993 -807 5969
rect -773 4993 -761 5969
rect -819 4981 -761 4993
rect -661 5969 -603 5981
rect -661 4993 -649 5969
rect -615 4993 -603 5969
rect -661 4981 -603 4993
rect -503 5969 -445 5981
rect -503 4993 -491 5969
rect -457 4993 -445 5969
rect -503 4981 -445 4993
rect -345 5969 -287 5981
rect -345 4993 -333 5969
rect -299 4993 -287 5969
rect -345 4981 -287 4993
rect -187 5969 -129 5981
rect -187 4993 -175 5969
rect -141 4993 -129 5969
rect -187 4981 -129 4993
rect -29 5969 29 5981
rect -29 4993 -17 5969
rect 17 4993 29 5969
rect -29 4981 29 4993
rect 129 5969 187 5981
rect 129 4993 141 5969
rect 175 4993 187 5969
rect 129 4981 187 4993
rect 287 5969 345 5981
rect 287 4993 299 5969
rect 333 4993 345 5969
rect 287 4981 345 4993
rect 445 5969 503 5981
rect 445 4993 457 5969
rect 491 4993 503 5969
rect 445 4981 503 4993
rect 603 5969 661 5981
rect 603 4993 615 5969
rect 649 4993 661 5969
rect 603 4981 661 4993
rect 761 5969 819 5981
rect 761 4993 773 5969
rect 807 4993 819 5969
rect 761 4981 819 4993
rect 919 5969 977 5981
rect 919 4993 931 5969
rect 965 4993 977 5969
rect 919 4981 977 4993
rect 1077 5969 1135 5981
rect 1077 4993 1089 5969
rect 1123 4993 1135 5969
rect 1077 4981 1135 4993
rect 1235 5969 1293 5981
rect 1235 4993 1247 5969
rect 1281 4993 1293 5969
rect 1235 4981 1293 4993
rect 1393 5969 1451 5981
rect 1393 4993 1405 5969
rect 1439 4993 1451 5969
rect 1393 4981 1451 4993
rect 1551 5969 1609 5981
rect 1551 4993 1563 5969
rect 1597 4993 1609 5969
rect 1551 4981 1609 4993
rect -1609 4751 -1551 4763
rect -1609 3775 -1597 4751
rect -1563 3775 -1551 4751
rect -1609 3763 -1551 3775
rect -1451 4751 -1393 4763
rect -1451 3775 -1439 4751
rect -1405 3775 -1393 4751
rect -1451 3763 -1393 3775
rect -1293 4751 -1235 4763
rect -1293 3775 -1281 4751
rect -1247 3775 -1235 4751
rect -1293 3763 -1235 3775
rect -1135 4751 -1077 4763
rect -1135 3775 -1123 4751
rect -1089 3775 -1077 4751
rect -1135 3763 -1077 3775
rect -977 4751 -919 4763
rect -977 3775 -965 4751
rect -931 3775 -919 4751
rect -977 3763 -919 3775
rect -819 4751 -761 4763
rect -819 3775 -807 4751
rect -773 3775 -761 4751
rect -819 3763 -761 3775
rect -661 4751 -603 4763
rect -661 3775 -649 4751
rect -615 3775 -603 4751
rect -661 3763 -603 3775
rect -503 4751 -445 4763
rect -503 3775 -491 4751
rect -457 3775 -445 4751
rect -503 3763 -445 3775
rect -345 4751 -287 4763
rect -345 3775 -333 4751
rect -299 3775 -287 4751
rect -345 3763 -287 3775
rect -187 4751 -129 4763
rect -187 3775 -175 4751
rect -141 3775 -129 4751
rect -187 3763 -129 3775
rect -29 4751 29 4763
rect -29 3775 -17 4751
rect 17 3775 29 4751
rect -29 3763 29 3775
rect 129 4751 187 4763
rect 129 3775 141 4751
rect 175 3775 187 4751
rect 129 3763 187 3775
rect 287 4751 345 4763
rect 287 3775 299 4751
rect 333 3775 345 4751
rect 287 3763 345 3775
rect 445 4751 503 4763
rect 445 3775 457 4751
rect 491 3775 503 4751
rect 445 3763 503 3775
rect 603 4751 661 4763
rect 603 3775 615 4751
rect 649 3775 661 4751
rect 603 3763 661 3775
rect 761 4751 819 4763
rect 761 3775 773 4751
rect 807 3775 819 4751
rect 761 3763 819 3775
rect 919 4751 977 4763
rect 919 3775 931 4751
rect 965 3775 977 4751
rect 919 3763 977 3775
rect 1077 4751 1135 4763
rect 1077 3775 1089 4751
rect 1123 3775 1135 4751
rect 1077 3763 1135 3775
rect 1235 4751 1293 4763
rect 1235 3775 1247 4751
rect 1281 3775 1293 4751
rect 1235 3763 1293 3775
rect 1393 4751 1451 4763
rect 1393 3775 1405 4751
rect 1439 3775 1451 4751
rect 1393 3763 1451 3775
rect 1551 4751 1609 4763
rect 1551 3775 1563 4751
rect 1597 3775 1609 4751
rect 1551 3763 1609 3775
rect -1609 3533 -1551 3545
rect -1609 2557 -1597 3533
rect -1563 2557 -1551 3533
rect -1609 2545 -1551 2557
rect -1451 3533 -1393 3545
rect -1451 2557 -1439 3533
rect -1405 2557 -1393 3533
rect -1451 2545 -1393 2557
rect -1293 3533 -1235 3545
rect -1293 2557 -1281 3533
rect -1247 2557 -1235 3533
rect -1293 2545 -1235 2557
rect -1135 3533 -1077 3545
rect -1135 2557 -1123 3533
rect -1089 2557 -1077 3533
rect -1135 2545 -1077 2557
rect -977 3533 -919 3545
rect -977 2557 -965 3533
rect -931 2557 -919 3533
rect -977 2545 -919 2557
rect -819 3533 -761 3545
rect -819 2557 -807 3533
rect -773 2557 -761 3533
rect -819 2545 -761 2557
rect -661 3533 -603 3545
rect -661 2557 -649 3533
rect -615 2557 -603 3533
rect -661 2545 -603 2557
rect -503 3533 -445 3545
rect -503 2557 -491 3533
rect -457 2557 -445 3533
rect -503 2545 -445 2557
rect -345 3533 -287 3545
rect -345 2557 -333 3533
rect -299 2557 -287 3533
rect -345 2545 -287 2557
rect -187 3533 -129 3545
rect -187 2557 -175 3533
rect -141 2557 -129 3533
rect -187 2545 -129 2557
rect -29 3533 29 3545
rect -29 2557 -17 3533
rect 17 2557 29 3533
rect -29 2545 29 2557
rect 129 3533 187 3545
rect 129 2557 141 3533
rect 175 2557 187 3533
rect 129 2545 187 2557
rect 287 3533 345 3545
rect 287 2557 299 3533
rect 333 2557 345 3533
rect 287 2545 345 2557
rect 445 3533 503 3545
rect 445 2557 457 3533
rect 491 2557 503 3533
rect 445 2545 503 2557
rect 603 3533 661 3545
rect 603 2557 615 3533
rect 649 2557 661 3533
rect 603 2545 661 2557
rect 761 3533 819 3545
rect 761 2557 773 3533
rect 807 2557 819 3533
rect 761 2545 819 2557
rect 919 3533 977 3545
rect 919 2557 931 3533
rect 965 2557 977 3533
rect 919 2545 977 2557
rect 1077 3533 1135 3545
rect 1077 2557 1089 3533
rect 1123 2557 1135 3533
rect 1077 2545 1135 2557
rect 1235 3533 1293 3545
rect 1235 2557 1247 3533
rect 1281 2557 1293 3533
rect 1235 2545 1293 2557
rect 1393 3533 1451 3545
rect 1393 2557 1405 3533
rect 1439 2557 1451 3533
rect 1393 2545 1451 2557
rect 1551 3533 1609 3545
rect 1551 2557 1563 3533
rect 1597 2557 1609 3533
rect 1551 2545 1609 2557
rect -1609 2315 -1551 2327
rect -1609 1339 -1597 2315
rect -1563 1339 -1551 2315
rect -1609 1327 -1551 1339
rect -1451 2315 -1393 2327
rect -1451 1339 -1439 2315
rect -1405 1339 -1393 2315
rect -1451 1327 -1393 1339
rect -1293 2315 -1235 2327
rect -1293 1339 -1281 2315
rect -1247 1339 -1235 2315
rect -1293 1327 -1235 1339
rect -1135 2315 -1077 2327
rect -1135 1339 -1123 2315
rect -1089 1339 -1077 2315
rect -1135 1327 -1077 1339
rect -977 2315 -919 2327
rect -977 1339 -965 2315
rect -931 1339 -919 2315
rect -977 1327 -919 1339
rect -819 2315 -761 2327
rect -819 1339 -807 2315
rect -773 1339 -761 2315
rect -819 1327 -761 1339
rect -661 2315 -603 2327
rect -661 1339 -649 2315
rect -615 1339 -603 2315
rect -661 1327 -603 1339
rect -503 2315 -445 2327
rect -503 1339 -491 2315
rect -457 1339 -445 2315
rect -503 1327 -445 1339
rect -345 2315 -287 2327
rect -345 1339 -333 2315
rect -299 1339 -287 2315
rect -345 1327 -287 1339
rect -187 2315 -129 2327
rect -187 1339 -175 2315
rect -141 1339 -129 2315
rect -187 1327 -129 1339
rect -29 2315 29 2327
rect -29 1339 -17 2315
rect 17 1339 29 2315
rect -29 1327 29 1339
rect 129 2315 187 2327
rect 129 1339 141 2315
rect 175 1339 187 2315
rect 129 1327 187 1339
rect 287 2315 345 2327
rect 287 1339 299 2315
rect 333 1339 345 2315
rect 287 1327 345 1339
rect 445 2315 503 2327
rect 445 1339 457 2315
rect 491 1339 503 2315
rect 445 1327 503 1339
rect 603 2315 661 2327
rect 603 1339 615 2315
rect 649 1339 661 2315
rect 603 1327 661 1339
rect 761 2315 819 2327
rect 761 1339 773 2315
rect 807 1339 819 2315
rect 761 1327 819 1339
rect 919 2315 977 2327
rect 919 1339 931 2315
rect 965 1339 977 2315
rect 919 1327 977 1339
rect 1077 2315 1135 2327
rect 1077 1339 1089 2315
rect 1123 1339 1135 2315
rect 1077 1327 1135 1339
rect 1235 2315 1293 2327
rect 1235 1339 1247 2315
rect 1281 1339 1293 2315
rect 1235 1327 1293 1339
rect 1393 2315 1451 2327
rect 1393 1339 1405 2315
rect 1439 1339 1451 2315
rect 1393 1327 1451 1339
rect 1551 2315 1609 2327
rect 1551 1339 1563 2315
rect 1597 1339 1609 2315
rect 1551 1327 1609 1339
rect -1609 1097 -1551 1109
rect -1609 121 -1597 1097
rect -1563 121 -1551 1097
rect -1609 109 -1551 121
rect -1451 1097 -1393 1109
rect -1451 121 -1439 1097
rect -1405 121 -1393 1097
rect -1451 109 -1393 121
rect -1293 1097 -1235 1109
rect -1293 121 -1281 1097
rect -1247 121 -1235 1097
rect -1293 109 -1235 121
rect -1135 1097 -1077 1109
rect -1135 121 -1123 1097
rect -1089 121 -1077 1097
rect -1135 109 -1077 121
rect -977 1097 -919 1109
rect -977 121 -965 1097
rect -931 121 -919 1097
rect -977 109 -919 121
rect -819 1097 -761 1109
rect -819 121 -807 1097
rect -773 121 -761 1097
rect -819 109 -761 121
rect -661 1097 -603 1109
rect -661 121 -649 1097
rect -615 121 -603 1097
rect -661 109 -603 121
rect -503 1097 -445 1109
rect -503 121 -491 1097
rect -457 121 -445 1097
rect -503 109 -445 121
rect -345 1097 -287 1109
rect -345 121 -333 1097
rect -299 121 -287 1097
rect -345 109 -287 121
rect -187 1097 -129 1109
rect -187 121 -175 1097
rect -141 121 -129 1097
rect -187 109 -129 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 129 1097 187 1109
rect 129 121 141 1097
rect 175 121 187 1097
rect 129 109 187 121
rect 287 1097 345 1109
rect 287 121 299 1097
rect 333 121 345 1097
rect 287 109 345 121
rect 445 1097 503 1109
rect 445 121 457 1097
rect 491 121 503 1097
rect 445 109 503 121
rect 603 1097 661 1109
rect 603 121 615 1097
rect 649 121 661 1097
rect 603 109 661 121
rect 761 1097 819 1109
rect 761 121 773 1097
rect 807 121 819 1097
rect 761 109 819 121
rect 919 1097 977 1109
rect 919 121 931 1097
rect 965 121 977 1097
rect 919 109 977 121
rect 1077 1097 1135 1109
rect 1077 121 1089 1097
rect 1123 121 1135 1097
rect 1077 109 1135 121
rect 1235 1097 1293 1109
rect 1235 121 1247 1097
rect 1281 121 1293 1097
rect 1235 109 1293 121
rect 1393 1097 1451 1109
rect 1393 121 1405 1097
rect 1439 121 1451 1097
rect 1393 109 1451 121
rect 1551 1097 1609 1109
rect 1551 121 1563 1097
rect 1597 121 1609 1097
rect 1551 109 1609 121
rect -1609 -121 -1551 -109
rect -1609 -1097 -1597 -121
rect -1563 -1097 -1551 -121
rect -1609 -1109 -1551 -1097
rect -1451 -121 -1393 -109
rect -1451 -1097 -1439 -121
rect -1405 -1097 -1393 -121
rect -1451 -1109 -1393 -1097
rect -1293 -121 -1235 -109
rect -1293 -1097 -1281 -121
rect -1247 -1097 -1235 -121
rect -1293 -1109 -1235 -1097
rect -1135 -121 -1077 -109
rect -1135 -1097 -1123 -121
rect -1089 -1097 -1077 -121
rect -1135 -1109 -1077 -1097
rect -977 -121 -919 -109
rect -977 -1097 -965 -121
rect -931 -1097 -919 -121
rect -977 -1109 -919 -1097
rect -819 -121 -761 -109
rect -819 -1097 -807 -121
rect -773 -1097 -761 -121
rect -819 -1109 -761 -1097
rect -661 -121 -603 -109
rect -661 -1097 -649 -121
rect -615 -1097 -603 -121
rect -661 -1109 -603 -1097
rect -503 -121 -445 -109
rect -503 -1097 -491 -121
rect -457 -1097 -445 -121
rect -503 -1109 -445 -1097
rect -345 -121 -287 -109
rect -345 -1097 -333 -121
rect -299 -1097 -287 -121
rect -345 -1109 -287 -1097
rect -187 -121 -129 -109
rect -187 -1097 -175 -121
rect -141 -1097 -129 -121
rect -187 -1109 -129 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 129 -121 187 -109
rect 129 -1097 141 -121
rect 175 -1097 187 -121
rect 129 -1109 187 -1097
rect 287 -121 345 -109
rect 287 -1097 299 -121
rect 333 -1097 345 -121
rect 287 -1109 345 -1097
rect 445 -121 503 -109
rect 445 -1097 457 -121
rect 491 -1097 503 -121
rect 445 -1109 503 -1097
rect 603 -121 661 -109
rect 603 -1097 615 -121
rect 649 -1097 661 -121
rect 603 -1109 661 -1097
rect 761 -121 819 -109
rect 761 -1097 773 -121
rect 807 -1097 819 -121
rect 761 -1109 819 -1097
rect 919 -121 977 -109
rect 919 -1097 931 -121
rect 965 -1097 977 -121
rect 919 -1109 977 -1097
rect 1077 -121 1135 -109
rect 1077 -1097 1089 -121
rect 1123 -1097 1135 -121
rect 1077 -1109 1135 -1097
rect 1235 -121 1293 -109
rect 1235 -1097 1247 -121
rect 1281 -1097 1293 -121
rect 1235 -1109 1293 -1097
rect 1393 -121 1451 -109
rect 1393 -1097 1405 -121
rect 1439 -1097 1451 -121
rect 1393 -1109 1451 -1097
rect 1551 -121 1609 -109
rect 1551 -1097 1563 -121
rect 1597 -1097 1609 -121
rect 1551 -1109 1609 -1097
rect -1609 -1339 -1551 -1327
rect -1609 -2315 -1597 -1339
rect -1563 -2315 -1551 -1339
rect -1609 -2327 -1551 -2315
rect -1451 -1339 -1393 -1327
rect -1451 -2315 -1439 -1339
rect -1405 -2315 -1393 -1339
rect -1451 -2327 -1393 -2315
rect -1293 -1339 -1235 -1327
rect -1293 -2315 -1281 -1339
rect -1247 -2315 -1235 -1339
rect -1293 -2327 -1235 -2315
rect -1135 -1339 -1077 -1327
rect -1135 -2315 -1123 -1339
rect -1089 -2315 -1077 -1339
rect -1135 -2327 -1077 -2315
rect -977 -1339 -919 -1327
rect -977 -2315 -965 -1339
rect -931 -2315 -919 -1339
rect -977 -2327 -919 -2315
rect -819 -1339 -761 -1327
rect -819 -2315 -807 -1339
rect -773 -2315 -761 -1339
rect -819 -2327 -761 -2315
rect -661 -1339 -603 -1327
rect -661 -2315 -649 -1339
rect -615 -2315 -603 -1339
rect -661 -2327 -603 -2315
rect -503 -1339 -445 -1327
rect -503 -2315 -491 -1339
rect -457 -2315 -445 -1339
rect -503 -2327 -445 -2315
rect -345 -1339 -287 -1327
rect -345 -2315 -333 -1339
rect -299 -2315 -287 -1339
rect -345 -2327 -287 -2315
rect -187 -1339 -129 -1327
rect -187 -2315 -175 -1339
rect -141 -2315 -129 -1339
rect -187 -2327 -129 -2315
rect -29 -1339 29 -1327
rect -29 -2315 -17 -1339
rect 17 -2315 29 -1339
rect -29 -2327 29 -2315
rect 129 -1339 187 -1327
rect 129 -2315 141 -1339
rect 175 -2315 187 -1339
rect 129 -2327 187 -2315
rect 287 -1339 345 -1327
rect 287 -2315 299 -1339
rect 333 -2315 345 -1339
rect 287 -2327 345 -2315
rect 445 -1339 503 -1327
rect 445 -2315 457 -1339
rect 491 -2315 503 -1339
rect 445 -2327 503 -2315
rect 603 -1339 661 -1327
rect 603 -2315 615 -1339
rect 649 -2315 661 -1339
rect 603 -2327 661 -2315
rect 761 -1339 819 -1327
rect 761 -2315 773 -1339
rect 807 -2315 819 -1339
rect 761 -2327 819 -2315
rect 919 -1339 977 -1327
rect 919 -2315 931 -1339
rect 965 -2315 977 -1339
rect 919 -2327 977 -2315
rect 1077 -1339 1135 -1327
rect 1077 -2315 1089 -1339
rect 1123 -2315 1135 -1339
rect 1077 -2327 1135 -2315
rect 1235 -1339 1293 -1327
rect 1235 -2315 1247 -1339
rect 1281 -2315 1293 -1339
rect 1235 -2327 1293 -2315
rect 1393 -1339 1451 -1327
rect 1393 -2315 1405 -1339
rect 1439 -2315 1451 -1339
rect 1393 -2327 1451 -2315
rect 1551 -1339 1609 -1327
rect 1551 -2315 1563 -1339
rect 1597 -2315 1609 -1339
rect 1551 -2327 1609 -2315
rect -1609 -2557 -1551 -2545
rect -1609 -3533 -1597 -2557
rect -1563 -3533 -1551 -2557
rect -1609 -3545 -1551 -3533
rect -1451 -2557 -1393 -2545
rect -1451 -3533 -1439 -2557
rect -1405 -3533 -1393 -2557
rect -1451 -3545 -1393 -3533
rect -1293 -2557 -1235 -2545
rect -1293 -3533 -1281 -2557
rect -1247 -3533 -1235 -2557
rect -1293 -3545 -1235 -3533
rect -1135 -2557 -1077 -2545
rect -1135 -3533 -1123 -2557
rect -1089 -3533 -1077 -2557
rect -1135 -3545 -1077 -3533
rect -977 -2557 -919 -2545
rect -977 -3533 -965 -2557
rect -931 -3533 -919 -2557
rect -977 -3545 -919 -3533
rect -819 -2557 -761 -2545
rect -819 -3533 -807 -2557
rect -773 -3533 -761 -2557
rect -819 -3545 -761 -3533
rect -661 -2557 -603 -2545
rect -661 -3533 -649 -2557
rect -615 -3533 -603 -2557
rect -661 -3545 -603 -3533
rect -503 -2557 -445 -2545
rect -503 -3533 -491 -2557
rect -457 -3533 -445 -2557
rect -503 -3545 -445 -3533
rect -345 -2557 -287 -2545
rect -345 -3533 -333 -2557
rect -299 -3533 -287 -2557
rect -345 -3545 -287 -3533
rect -187 -2557 -129 -2545
rect -187 -3533 -175 -2557
rect -141 -3533 -129 -2557
rect -187 -3545 -129 -3533
rect -29 -2557 29 -2545
rect -29 -3533 -17 -2557
rect 17 -3533 29 -2557
rect -29 -3545 29 -3533
rect 129 -2557 187 -2545
rect 129 -3533 141 -2557
rect 175 -3533 187 -2557
rect 129 -3545 187 -3533
rect 287 -2557 345 -2545
rect 287 -3533 299 -2557
rect 333 -3533 345 -2557
rect 287 -3545 345 -3533
rect 445 -2557 503 -2545
rect 445 -3533 457 -2557
rect 491 -3533 503 -2557
rect 445 -3545 503 -3533
rect 603 -2557 661 -2545
rect 603 -3533 615 -2557
rect 649 -3533 661 -2557
rect 603 -3545 661 -3533
rect 761 -2557 819 -2545
rect 761 -3533 773 -2557
rect 807 -3533 819 -2557
rect 761 -3545 819 -3533
rect 919 -2557 977 -2545
rect 919 -3533 931 -2557
rect 965 -3533 977 -2557
rect 919 -3545 977 -3533
rect 1077 -2557 1135 -2545
rect 1077 -3533 1089 -2557
rect 1123 -3533 1135 -2557
rect 1077 -3545 1135 -3533
rect 1235 -2557 1293 -2545
rect 1235 -3533 1247 -2557
rect 1281 -3533 1293 -2557
rect 1235 -3545 1293 -3533
rect 1393 -2557 1451 -2545
rect 1393 -3533 1405 -2557
rect 1439 -3533 1451 -2557
rect 1393 -3545 1451 -3533
rect 1551 -2557 1609 -2545
rect 1551 -3533 1563 -2557
rect 1597 -3533 1609 -2557
rect 1551 -3545 1609 -3533
rect -1609 -3775 -1551 -3763
rect -1609 -4751 -1597 -3775
rect -1563 -4751 -1551 -3775
rect -1609 -4763 -1551 -4751
rect -1451 -3775 -1393 -3763
rect -1451 -4751 -1439 -3775
rect -1405 -4751 -1393 -3775
rect -1451 -4763 -1393 -4751
rect -1293 -3775 -1235 -3763
rect -1293 -4751 -1281 -3775
rect -1247 -4751 -1235 -3775
rect -1293 -4763 -1235 -4751
rect -1135 -3775 -1077 -3763
rect -1135 -4751 -1123 -3775
rect -1089 -4751 -1077 -3775
rect -1135 -4763 -1077 -4751
rect -977 -3775 -919 -3763
rect -977 -4751 -965 -3775
rect -931 -4751 -919 -3775
rect -977 -4763 -919 -4751
rect -819 -3775 -761 -3763
rect -819 -4751 -807 -3775
rect -773 -4751 -761 -3775
rect -819 -4763 -761 -4751
rect -661 -3775 -603 -3763
rect -661 -4751 -649 -3775
rect -615 -4751 -603 -3775
rect -661 -4763 -603 -4751
rect -503 -3775 -445 -3763
rect -503 -4751 -491 -3775
rect -457 -4751 -445 -3775
rect -503 -4763 -445 -4751
rect -345 -3775 -287 -3763
rect -345 -4751 -333 -3775
rect -299 -4751 -287 -3775
rect -345 -4763 -287 -4751
rect -187 -3775 -129 -3763
rect -187 -4751 -175 -3775
rect -141 -4751 -129 -3775
rect -187 -4763 -129 -4751
rect -29 -3775 29 -3763
rect -29 -4751 -17 -3775
rect 17 -4751 29 -3775
rect -29 -4763 29 -4751
rect 129 -3775 187 -3763
rect 129 -4751 141 -3775
rect 175 -4751 187 -3775
rect 129 -4763 187 -4751
rect 287 -3775 345 -3763
rect 287 -4751 299 -3775
rect 333 -4751 345 -3775
rect 287 -4763 345 -4751
rect 445 -3775 503 -3763
rect 445 -4751 457 -3775
rect 491 -4751 503 -3775
rect 445 -4763 503 -4751
rect 603 -3775 661 -3763
rect 603 -4751 615 -3775
rect 649 -4751 661 -3775
rect 603 -4763 661 -4751
rect 761 -3775 819 -3763
rect 761 -4751 773 -3775
rect 807 -4751 819 -3775
rect 761 -4763 819 -4751
rect 919 -3775 977 -3763
rect 919 -4751 931 -3775
rect 965 -4751 977 -3775
rect 919 -4763 977 -4751
rect 1077 -3775 1135 -3763
rect 1077 -4751 1089 -3775
rect 1123 -4751 1135 -3775
rect 1077 -4763 1135 -4751
rect 1235 -3775 1293 -3763
rect 1235 -4751 1247 -3775
rect 1281 -4751 1293 -3775
rect 1235 -4763 1293 -4751
rect 1393 -3775 1451 -3763
rect 1393 -4751 1405 -3775
rect 1439 -4751 1451 -3775
rect 1393 -4763 1451 -4751
rect 1551 -3775 1609 -3763
rect 1551 -4751 1563 -3775
rect 1597 -4751 1609 -3775
rect 1551 -4763 1609 -4751
rect -1609 -4993 -1551 -4981
rect -1609 -5969 -1597 -4993
rect -1563 -5969 -1551 -4993
rect -1609 -5981 -1551 -5969
rect -1451 -4993 -1393 -4981
rect -1451 -5969 -1439 -4993
rect -1405 -5969 -1393 -4993
rect -1451 -5981 -1393 -5969
rect -1293 -4993 -1235 -4981
rect -1293 -5969 -1281 -4993
rect -1247 -5969 -1235 -4993
rect -1293 -5981 -1235 -5969
rect -1135 -4993 -1077 -4981
rect -1135 -5969 -1123 -4993
rect -1089 -5969 -1077 -4993
rect -1135 -5981 -1077 -5969
rect -977 -4993 -919 -4981
rect -977 -5969 -965 -4993
rect -931 -5969 -919 -4993
rect -977 -5981 -919 -5969
rect -819 -4993 -761 -4981
rect -819 -5969 -807 -4993
rect -773 -5969 -761 -4993
rect -819 -5981 -761 -5969
rect -661 -4993 -603 -4981
rect -661 -5969 -649 -4993
rect -615 -5969 -603 -4993
rect -661 -5981 -603 -5969
rect -503 -4993 -445 -4981
rect -503 -5969 -491 -4993
rect -457 -5969 -445 -4993
rect -503 -5981 -445 -5969
rect -345 -4993 -287 -4981
rect -345 -5969 -333 -4993
rect -299 -5969 -287 -4993
rect -345 -5981 -287 -5969
rect -187 -4993 -129 -4981
rect -187 -5969 -175 -4993
rect -141 -5969 -129 -4993
rect -187 -5981 -129 -5969
rect -29 -4993 29 -4981
rect -29 -5969 -17 -4993
rect 17 -5969 29 -4993
rect -29 -5981 29 -5969
rect 129 -4993 187 -4981
rect 129 -5969 141 -4993
rect 175 -5969 187 -4993
rect 129 -5981 187 -5969
rect 287 -4993 345 -4981
rect 287 -5969 299 -4993
rect 333 -5969 345 -4993
rect 287 -5981 345 -5969
rect 445 -4993 503 -4981
rect 445 -5969 457 -4993
rect 491 -5969 503 -4993
rect 445 -5981 503 -5969
rect 603 -4993 661 -4981
rect 603 -5969 615 -4993
rect 649 -5969 661 -4993
rect 603 -5981 661 -5969
rect 761 -4993 819 -4981
rect 761 -5969 773 -4993
rect 807 -5969 819 -4993
rect 761 -5981 819 -5969
rect 919 -4993 977 -4981
rect 919 -5969 931 -4993
rect 965 -5969 977 -4993
rect 919 -5981 977 -5969
rect 1077 -4993 1135 -4981
rect 1077 -5969 1089 -4993
rect 1123 -5969 1135 -4993
rect 1077 -5981 1135 -5969
rect 1235 -4993 1293 -4981
rect 1235 -5969 1247 -4993
rect 1281 -5969 1293 -4993
rect 1235 -5981 1293 -5969
rect 1393 -4993 1451 -4981
rect 1393 -5969 1405 -4993
rect 1439 -5969 1451 -4993
rect 1393 -5981 1451 -5969
rect 1551 -4993 1609 -4981
rect 1551 -5969 1563 -4993
rect 1597 -5969 1609 -4993
rect 1551 -5981 1609 -5969
<< mvndiffc >>
rect -1597 4993 -1563 5969
rect -1439 4993 -1405 5969
rect -1281 4993 -1247 5969
rect -1123 4993 -1089 5969
rect -965 4993 -931 5969
rect -807 4993 -773 5969
rect -649 4993 -615 5969
rect -491 4993 -457 5969
rect -333 4993 -299 5969
rect -175 4993 -141 5969
rect -17 4993 17 5969
rect 141 4993 175 5969
rect 299 4993 333 5969
rect 457 4993 491 5969
rect 615 4993 649 5969
rect 773 4993 807 5969
rect 931 4993 965 5969
rect 1089 4993 1123 5969
rect 1247 4993 1281 5969
rect 1405 4993 1439 5969
rect 1563 4993 1597 5969
rect -1597 3775 -1563 4751
rect -1439 3775 -1405 4751
rect -1281 3775 -1247 4751
rect -1123 3775 -1089 4751
rect -965 3775 -931 4751
rect -807 3775 -773 4751
rect -649 3775 -615 4751
rect -491 3775 -457 4751
rect -333 3775 -299 4751
rect -175 3775 -141 4751
rect -17 3775 17 4751
rect 141 3775 175 4751
rect 299 3775 333 4751
rect 457 3775 491 4751
rect 615 3775 649 4751
rect 773 3775 807 4751
rect 931 3775 965 4751
rect 1089 3775 1123 4751
rect 1247 3775 1281 4751
rect 1405 3775 1439 4751
rect 1563 3775 1597 4751
rect -1597 2557 -1563 3533
rect -1439 2557 -1405 3533
rect -1281 2557 -1247 3533
rect -1123 2557 -1089 3533
rect -965 2557 -931 3533
rect -807 2557 -773 3533
rect -649 2557 -615 3533
rect -491 2557 -457 3533
rect -333 2557 -299 3533
rect -175 2557 -141 3533
rect -17 2557 17 3533
rect 141 2557 175 3533
rect 299 2557 333 3533
rect 457 2557 491 3533
rect 615 2557 649 3533
rect 773 2557 807 3533
rect 931 2557 965 3533
rect 1089 2557 1123 3533
rect 1247 2557 1281 3533
rect 1405 2557 1439 3533
rect 1563 2557 1597 3533
rect -1597 1339 -1563 2315
rect -1439 1339 -1405 2315
rect -1281 1339 -1247 2315
rect -1123 1339 -1089 2315
rect -965 1339 -931 2315
rect -807 1339 -773 2315
rect -649 1339 -615 2315
rect -491 1339 -457 2315
rect -333 1339 -299 2315
rect -175 1339 -141 2315
rect -17 1339 17 2315
rect 141 1339 175 2315
rect 299 1339 333 2315
rect 457 1339 491 2315
rect 615 1339 649 2315
rect 773 1339 807 2315
rect 931 1339 965 2315
rect 1089 1339 1123 2315
rect 1247 1339 1281 2315
rect 1405 1339 1439 2315
rect 1563 1339 1597 2315
rect -1597 121 -1563 1097
rect -1439 121 -1405 1097
rect -1281 121 -1247 1097
rect -1123 121 -1089 1097
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect 1089 121 1123 1097
rect 1247 121 1281 1097
rect 1405 121 1439 1097
rect 1563 121 1597 1097
rect -1597 -1097 -1563 -121
rect -1439 -1097 -1405 -121
rect -1281 -1097 -1247 -121
rect -1123 -1097 -1089 -121
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
rect 1089 -1097 1123 -121
rect 1247 -1097 1281 -121
rect 1405 -1097 1439 -121
rect 1563 -1097 1597 -121
rect -1597 -2315 -1563 -1339
rect -1439 -2315 -1405 -1339
rect -1281 -2315 -1247 -1339
rect -1123 -2315 -1089 -1339
rect -965 -2315 -931 -1339
rect -807 -2315 -773 -1339
rect -649 -2315 -615 -1339
rect -491 -2315 -457 -1339
rect -333 -2315 -299 -1339
rect -175 -2315 -141 -1339
rect -17 -2315 17 -1339
rect 141 -2315 175 -1339
rect 299 -2315 333 -1339
rect 457 -2315 491 -1339
rect 615 -2315 649 -1339
rect 773 -2315 807 -1339
rect 931 -2315 965 -1339
rect 1089 -2315 1123 -1339
rect 1247 -2315 1281 -1339
rect 1405 -2315 1439 -1339
rect 1563 -2315 1597 -1339
rect -1597 -3533 -1563 -2557
rect -1439 -3533 -1405 -2557
rect -1281 -3533 -1247 -2557
rect -1123 -3533 -1089 -2557
rect -965 -3533 -931 -2557
rect -807 -3533 -773 -2557
rect -649 -3533 -615 -2557
rect -491 -3533 -457 -2557
rect -333 -3533 -299 -2557
rect -175 -3533 -141 -2557
rect -17 -3533 17 -2557
rect 141 -3533 175 -2557
rect 299 -3533 333 -2557
rect 457 -3533 491 -2557
rect 615 -3533 649 -2557
rect 773 -3533 807 -2557
rect 931 -3533 965 -2557
rect 1089 -3533 1123 -2557
rect 1247 -3533 1281 -2557
rect 1405 -3533 1439 -2557
rect 1563 -3533 1597 -2557
rect -1597 -4751 -1563 -3775
rect -1439 -4751 -1405 -3775
rect -1281 -4751 -1247 -3775
rect -1123 -4751 -1089 -3775
rect -965 -4751 -931 -3775
rect -807 -4751 -773 -3775
rect -649 -4751 -615 -3775
rect -491 -4751 -457 -3775
rect -333 -4751 -299 -3775
rect -175 -4751 -141 -3775
rect -17 -4751 17 -3775
rect 141 -4751 175 -3775
rect 299 -4751 333 -3775
rect 457 -4751 491 -3775
rect 615 -4751 649 -3775
rect 773 -4751 807 -3775
rect 931 -4751 965 -3775
rect 1089 -4751 1123 -3775
rect 1247 -4751 1281 -3775
rect 1405 -4751 1439 -3775
rect 1563 -4751 1597 -3775
rect -1597 -5969 -1563 -4993
rect -1439 -5969 -1405 -4993
rect -1281 -5969 -1247 -4993
rect -1123 -5969 -1089 -4993
rect -965 -5969 -931 -4993
rect -807 -5969 -773 -4993
rect -649 -5969 -615 -4993
rect -491 -5969 -457 -4993
rect -333 -5969 -299 -4993
rect -175 -5969 -141 -4993
rect -17 -5969 17 -4993
rect 141 -5969 175 -4993
rect 299 -5969 333 -4993
rect 457 -5969 491 -4993
rect 615 -5969 649 -4993
rect 773 -5969 807 -4993
rect 931 -5969 965 -4993
rect 1089 -5969 1123 -4993
rect 1247 -5969 1281 -4993
rect 1405 -5969 1439 -4993
rect 1563 -5969 1597 -4993
<< mvpsubdiff >>
rect -1753 6191 1753 6203
rect -1753 6157 -1645 6191
rect 1645 6157 1753 6191
rect -1753 6145 1753 6157
rect -1753 6095 -1695 6145
rect -1753 -6095 -1741 6095
rect -1707 -6095 -1695 6095
rect 1695 6095 1753 6145
rect -1753 -6145 -1695 -6095
rect 1695 -6095 1707 6095
rect 1741 -6095 1753 6095
rect 1695 -6145 1753 -6095
rect -1753 -6157 1753 -6145
rect -1753 -6191 -1645 -6157
rect 1645 -6191 1753 -6157
rect -1753 -6203 1753 -6191
<< mvpsubdiffcont >>
rect -1645 6157 1645 6191
rect -1741 -6095 -1707 6095
rect 1707 -6095 1741 6095
rect -1645 -6191 1645 -6157
<< poly >>
rect -1551 6053 -1451 6069
rect -1551 6019 -1535 6053
rect -1467 6019 -1451 6053
rect -1551 5981 -1451 6019
rect -1393 6053 -1293 6069
rect -1393 6019 -1377 6053
rect -1309 6019 -1293 6053
rect -1393 5981 -1293 6019
rect -1235 6053 -1135 6069
rect -1235 6019 -1219 6053
rect -1151 6019 -1135 6053
rect -1235 5981 -1135 6019
rect -1077 6053 -977 6069
rect -1077 6019 -1061 6053
rect -993 6019 -977 6053
rect -1077 5981 -977 6019
rect -919 6053 -819 6069
rect -919 6019 -903 6053
rect -835 6019 -819 6053
rect -919 5981 -819 6019
rect -761 6053 -661 6069
rect -761 6019 -745 6053
rect -677 6019 -661 6053
rect -761 5981 -661 6019
rect -603 6053 -503 6069
rect -603 6019 -587 6053
rect -519 6019 -503 6053
rect -603 5981 -503 6019
rect -445 6053 -345 6069
rect -445 6019 -429 6053
rect -361 6019 -345 6053
rect -445 5981 -345 6019
rect -287 6053 -187 6069
rect -287 6019 -271 6053
rect -203 6019 -187 6053
rect -287 5981 -187 6019
rect -129 6053 -29 6069
rect -129 6019 -113 6053
rect -45 6019 -29 6053
rect -129 5981 -29 6019
rect 29 6053 129 6069
rect 29 6019 45 6053
rect 113 6019 129 6053
rect 29 5981 129 6019
rect 187 6053 287 6069
rect 187 6019 203 6053
rect 271 6019 287 6053
rect 187 5981 287 6019
rect 345 6053 445 6069
rect 345 6019 361 6053
rect 429 6019 445 6053
rect 345 5981 445 6019
rect 503 6053 603 6069
rect 503 6019 519 6053
rect 587 6019 603 6053
rect 503 5981 603 6019
rect 661 6053 761 6069
rect 661 6019 677 6053
rect 745 6019 761 6053
rect 661 5981 761 6019
rect 819 6053 919 6069
rect 819 6019 835 6053
rect 903 6019 919 6053
rect 819 5981 919 6019
rect 977 6053 1077 6069
rect 977 6019 993 6053
rect 1061 6019 1077 6053
rect 977 5981 1077 6019
rect 1135 6053 1235 6069
rect 1135 6019 1151 6053
rect 1219 6019 1235 6053
rect 1135 5981 1235 6019
rect 1293 6053 1393 6069
rect 1293 6019 1309 6053
rect 1377 6019 1393 6053
rect 1293 5981 1393 6019
rect 1451 6053 1551 6069
rect 1451 6019 1467 6053
rect 1535 6019 1551 6053
rect 1451 5981 1551 6019
rect -1551 4943 -1451 4981
rect -1551 4909 -1535 4943
rect -1467 4909 -1451 4943
rect -1551 4893 -1451 4909
rect -1393 4943 -1293 4981
rect -1393 4909 -1377 4943
rect -1309 4909 -1293 4943
rect -1393 4893 -1293 4909
rect -1235 4943 -1135 4981
rect -1235 4909 -1219 4943
rect -1151 4909 -1135 4943
rect -1235 4893 -1135 4909
rect -1077 4943 -977 4981
rect -1077 4909 -1061 4943
rect -993 4909 -977 4943
rect -1077 4893 -977 4909
rect -919 4943 -819 4981
rect -919 4909 -903 4943
rect -835 4909 -819 4943
rect -919 4893 -819 4909
rect -761 4943 -661 4981
rect -761 4909 -745 4943
rect -677 4909 -661 4943
rect -761 4893 -661 4909
rect -603 4943 -503 4981
rect -603 4909 -587 4943
rect -519 4909 -503 4943
rect -603 4893 -503 4909
rect -445 4943 -345 4981
rect -445 4909 -429 4943
rect -361 4909 -345 4943
rect -445 4893 -345 4909
rect -287 4943 -187 4981
rect -287 4909 -271 4943
rect -203 4909 -187 4943
rect -287 4893 -187 4909
rect -129 4943 -29 4981
rect -129 4909 -113 4943
rect -45 4909 -29 4943
rect -129 4893 -29 4909
rect 29 4943 129 4981
rect 29 4909 45 4943
rect 113 4909 129 4943
rect 29 4893 129 4909
rect 187 4943 287 4981
rect 187 4909 203 4943
rect 271 4909 287 4943
rect 187 4893 287 4909
rect 345 4943 445 4981
rect 345 4909 361 4943
rect 429 4909 445 4943
rect 345 4893 445 4909
rect 503 4943 603 4981
rect 503 4909 519 4943
rect 587 4909 603 4943
rect 503 4893 603 4909
rect 661 4943 761 4981
rect 661 4909 677 4943
rect 745 4909 761 4943
rect 661 4893 761 4909
rect 819 4943 919 4981
rect 819 4909 835 4943
rect 903 4909 919 4943
rect 819 4893 919 4909
rect 977 4943 1077 4981
rect 977 4909 993 4943
rect 1061 4909 1077 4943
rect 977 4893 1077 4909
rect 1135 4943 1235 4981
rect 1135 4909 1151 4943
rect 1219 4909 1235 4943
rect 1135 4893 1235 4909
rect 1293 4943 1393 4981
rect 1293 4909 1309 4943
rect 1377 4909 1393 4943
rect 1293 4893 1393 4909
rect 1451 4943 1551 4981
rect 1451 4909 1467 4943
rect 1535 4909 1551 4943
rect 1451 4893 1551 4909
rect -1551 4835 -1451 4851
rect -1551 4801 -1535 4835
rect -1467 4801 -1451 4835
rect -1551 4763 -1451 4801
rect -1393 4835 -1293 4851
rect -1393 4801 -1377 4835
rect -1309 4801 -1293 4835
rect -1393 4763 -1293 4801
rect -1235 4835 -1135 4851
rect -1235 4801 -1219 4835
rect -1151 4801 -1135 4835
rect -1235 4763 -1135 4801
rect -1077 4835 -977 4851
rect -1077 4801 -1061 4835
rect -993 4801 -977 4835
rect -1077 4763 -977 4801
rect -919 4835 -819 4851
rect -919 4801 -903 4835
rect -835 4801 -819 4835
rect -919 4763 -819 4801
rect -761 4835 -661 4851
rect -761 4801 -745 4835
rect -677 4801 -661 4835
rect -761 4763 -661 4801
rect -603 4835 -503 4851
rect -603 4801 -587 4835
rect -519 4801 -503 4835
rect -603 4763 -503 4801
rect -445 4835 -345 4851
rect -445 4801 -429 4835
rect -361 4801 -345 4835
rect -445 4763 -345 4801
rect -287 4835 -187 4851
rect -287 4801 -271 4835
rect -203 4801 -187 4835
rect -287 4763 -187 4801
rect -129 4835 -29 4851
rect -129 4801 -113 4835
rect -45 4801 -29 4835
rect -129 4763 -29 4801
rect 29 4835 129 4851
rect 29 4801 45 4835
rect 113 4801 129 4835
rect 29 4763 129 4801
rect 187 4835 287 4851
rect 187 4801 203 4835
rect 271 4801 287 4835
rect 187 4763 287 4801
rect 345 4835 445 4851
rect 345 4801 361 4835
rect 429 4801 445 4835
rect 345 4763 445 4801
rect 503 4835 603 4851
rect 503 4801 519 4835
rect 587 4801 603 4835
rect 503 4763 603 4801
rect 661 4835 761 4851
rect 661 4801 677 4835
rect 745 4801 761 4835
rect 661 4763 761 4801
rect 819 4835 919 4851
rect 819 4801 835 4835
rect 903 4801 919 4835
rect 819 4763 919 4801
rect 977 4835 1077 4851
rect 977 4801 993 4835
rect 1061 4801 1077 4835
rect 977 4763 1077 4801
rect 1135 4835 1235 4851
rect 1135 4801 1151 4835
rect 1219 4801 1235 4835
rect 1135 4763 1235 4801
rect 1293 4835 1393 4851
rect 1293 4801 1309 4835
rect 1377 4801 1393 4835
rect 1293 4763 1393 4801
rect 1451 4835 1551 4851
rect 1451 4801 1467 4835
rect 1535 4801 1551 4835
rect 1451 4763 1551 4801
rect -1551 3725 -1451 3763
rect -1551 3691 -1535 3725
rect -1467 3691 -1451 3725
rect -1551 3675 -1451 3691
rect -1393 3725 -1293 3763
rect -1393 3691 -1377 3725
rect -1309 3691 -1293 3725
rect -1393 3675 -1293 3691
rect -1235 3725 -1135 3763
rect -1235 3691 -1219 3725
rect -1151 3691 -1135 3725
rect -1235 3675 -1135 3691
rect -1077 3725 -977 3763
rect -1077 3691 -1061 3725
rect -993 3691 -977 3725
rect -1077 3675 -977 3691
rect -919 3725 -819 3763
rect -919 3691 -903 3725
rect -835 3691 -819 3725
rect -919 3675 -819 3691
rect -761 3725 -661 3763
rect -761 3691 -745 3725
rect -677 3691 -661 3725
rect -761 3675 -661 3691
rect -603 3725 -503 3763
rect -603 3691 -587 3725
rect -519 3691 -503 3725
rect -603 3675 -503 3691
rect -445 3725 -345 3763
rect -445 3691 -429 3725
rect -361 3691 -345 3725
rect -445 3675 -345 3691
rect -287 3725 -187 3763
rect -287 3691 -271 3725
rect -203 3691 -187 3725
rect -287 3675 -187 3691
rect -129 3725 -29 3763
rect -129 3691 -113 3725
rect -45 3691 -29 3725
rect -129 3675 -29 3691
rect 29 3725 129 3763
rect 29 3691 45 3725
rect 113 3691 129 3725
rect 29 3675 129 3691
rect 187 3725 287 3763
rect 187 3691 203 3725
rect 271 3691 287 3725
rect 187 3675 287 3691
rect 345 3725 445 3763
rect 345 3691 361 3725
rect 429 3691 445 3725
rect 345 3675 445 3691
rect 503 3725 603 3763
rect 503 3691 519 3725
rect 587 3691 603 3725
rect 503 3675 603 3691
rect 661 3725 761 3763
rect 661 3691 677 3725
rect 745 3691 761 3725
rect 661 3675 761 3691
rect 819 3725 919 3763
rect 819 3691 835 3725
rect 903 3691 919 3725
rect 819 3675 919 3691
rect 977 3725 1077 3763
rect 977 3691 993 3725
rect 1061 3691 1077 3725
rect 977 3675 1077 3691
rect 1135 3725 1235 3763
rect 1135 3691 1151 3725
rect 1219 3691 1235 3725
rect 1135 3675 1235 3691
rect 1293 3725 1393 3763
rect 1293 3691 1309 3725
rect 1377 3691 1393 3725
rect 1293 3675 1393 3691
rect 1451 3725 1551 3763
rect 1451 3691 1467 3725
rect 1535 3691 1551 3725
rect 1451 3675 1551 3691
rect -1551 3617 -1451 3633
rect -1551 3583 -1535 3617
rect -1467 3583 -1451 3617
rect -1551 3545 -1451 3583
rect -1393 3617 -1293 3633
rect -1393 3583 -1377 3617
rect -1309 3583 -1293 3617
rect -1393 3545 -1293 3583
rect -1235 3617 -1135 3633
rect -1235 3583 -1219 3617
rect -1151 3583 -1135 3617
rect -1235 3545 -1135 3583
rect -1077 3617 -977 3633
rect -1077 3583 -1061 3617
rect -993 3583 -977 3617
rect -1077 3545 -977 3583
rect -919 3617 -819 3633
rect -919 3583 -903 3617
rect -835 3583 -819 3617
rect -919 3545 -819 3583
rect -761 3617 -661 3633
rect -761 3583 -745 3617
rect -677 3583 -661 3617
rect -761 3545 -661 3583
rect -603 3617 -503 3633
rect -603 3583 -587 3617
rect -519 3583 -503 3617
rect -603 3545 -503 3583
rect -445 3617 -345 3633
rect -445 3583 -429 3617
rect -361 3583 -345 3617
rect -445 3545 -345 3583
rect -287 3617 -187 3633
rect -287 3583 -271 3617
rect -203 3583 -187 3617
rect -287 3545 -187 3583
rect -129 3617 -29 3633
rect -129 3583 -113 3617
rect -45 3583 -29 3617
rect -129 3545 -29 3583
rect 29 3617 129 3633
rect 29 3583 45 3617
rect 113 3583 129 3617
rect 29 3545 129 3583
rect 187 3617 287 3633
rect 187 3583 203 3617
rect 271 3583 287 3617
rect 187 3545 287 3583
rect 345 3617 445 3633
rect 345 3583 361 3617
rect 429 3583 445 3617
rect 345 3545 445 3583
rect 503 3617 603 3633
rect 503 3583 519 3617
rect 587 3583 603 3617
rect 503 3545 603 3583
rect 661 3617 761 3633
rect 661 3583 677 3617
rect 745 3583 761 3617
rect 661 3545 761 3583
rect 819 3617 919 3633
rect 819 3583 835 3617
rect 903 3583 919 3617
rect 819 3545 919 3583
rect 977 3617 1077 3633
rect 977 3583 993 3617
rect 1061 3583 1077 3617
rect 977 3545 1077 3583
rect 1135 3617 1235 3633
rect 1135 3583 1151 3617
rect 1219 3583 1235 3617
rect 1135 3545 1235 3583
rect 1293 3617 1393 3633
rect 1293 3583 1309 3617
rect 1377 3583 1393 3617
rect 1293 3545 1393 3583
rect 1451 3617 1551 3633
rect 1451 3583 1467 3617
rect 1535 3583 1551 3617
rect 1451 3545 1551 3583
rect -1551 2507 -1451 2545
rect -1551 2473 -1535 2507
rect -1467 2473 -1451 2507
rect -1551 2457 -1451 2473
rect -1393 2507 -1293 2545
rect -1393 2473 -1377 2507
rect -1309 2473 -1293 2507
rect -1393 2457 -1293 2473
rect -1235 2507 -1135 2545
rect -1235 2473 -1219 2507
rect -1151 2473 -1135 2507
rect -1235 2457 -1135 2473
rect -1077 2507 -977 2545
rect -1077 2473 -1061 2507
rect -993 2473 -977 2507
rect -1077 2457 -977 2473
rect -919 2507 -819 2545
rect -919 2473 -903 2507
rect -835 2473 -819 2507
rect -919 2457 -819 2473
rect -761 2507 -661 2545
rect -761 2473 -745 2507
rect -677 2473 -661 2507
rect -761 2457 -661 2473
rect -603 2507 -503 2545
rect -603 2473 -587 2507
rect -519 2473 -503 2507
rect -603 2457 -503 2473
rect -445 2507 -345 2545
rect -445 2473 -429 2507
rect -361 2473 -345 2507
rect -445 2457 -345 2473
rect -287 2507 -187 2545
rect -287 2473 -271 2507
rect -203 2473 -187 2507
rect -287 2457 -187 2473
rect -129 2507 -29 2545
rect -129 2473 -113 2507
rect -45 2473 -29 2507
rect -129 2457 -29 2473
rect 29 2507 129 2545
rect 29 2473 45 2507
rect 113 2473 129 2507
rect 29 2457 129 2473
rect 187 2507 287 2545
rect 187 2473 203 2507
rect 271 2473 287 2507
rect 187 2457 287 2473
rect 345 2507 445 2545
rect 345 2473 361 2507
rect 429 2473 445 2507
rect 345 2457 445 2473
rect 503 2507 603 2545
rect 503 2473 519 2507
rect 587 2473 603 2507
rect 503 2457 603 2473
rect 661 2507 761 2545
rect 661 2473 677 2507
rect 745 2473 761 2507
rect 661 2457 761 2473
rect 819 2507 919 2545
rect 819 2473 835 2507
rect 903 2473 919 2507
rect 819 2457 919 2473
rect 977 2507 1077 2545
rect 977 2473 993 2507
rect 1061 2473 1077 2507
rect 977 2457 1077 2473
rect 1135 2507 1235 2545
rect 1135 2473 1151 2507
rect 1219 2473 1235 2507
rect 1135 2457 1235 2473
rect 1293 2507 1393 2545
rect 1293 2473 1309 2507
rect 1377 2473 1393 2507
rect 1293 2457 1393 2473
rect 1451 2507 1551 2545
rect 1451 2473 1467 2507
rect 1535 2473 1551 2507
rect 1451 2457 1551 2473
rect -1551 2399 -1451 2415
rect -1551 2365 -1535 2399
rect -1467 2365 -1451 2399
rect -1551 2327 -1451 2365
rect -1393 2399 -1293 2415
rect -1393 2365 -1377 2399
rect -1309 2365 -1293 2399
rect -1393 2327 -1293 2365
rect -1235 2399 -1135 2415
rect -1235 2365 -1219 2399
rect -1151 2365 -1135 2399
rect -1235 2327 -1135 2365
rect -1077 2399 -977 2415
rect -1077 2365 -1061 2399
rect -993 2365 -977 2399
rect -1077 2327 -977 2365
rect -919 2399 -819 2415
rect -919 2365 -903 2399
rect -835 2365 -819 2399
rect -919 2327 -819 2365
rect -761 2399 -661 2415
rect -761 2365 -745 2399
rect -677 2365 -661 2399
rect -761 2327 -661 2365
rect -603 2399 -503 2415
rect -603 2365 -587 2399
rect -519 2365 -503 2399
rect -603 2327 -503 2365
rect -445 2399 -345 2415
rect -445 2365 -429 2399
rect -361 2365 -345 2399
rect -445 2327 -345 2365
rect -287 2399 -187 2415
rect -287 2365 -271 2399
rect -203 2365 -187 2399
rect -287 2327 -187 2365
rect -129 2399 -29 2415
rect -129 2365 -113 2399
rect -45 2365 -29 2399
rect -129 2327 -29 2365
rect 29 2399 129 2415
rect 29 2365 45 2399
rect 113 2365 129 2399
rect 29 2327 129 2365
rect 187 2399 287 2415
rect 187 2365 203 2399
rect 271 2365 287 2399
rect 187 2327 287 2365
rect 345 2399 445 2415
rect 345 2365 361 2399
rect 429 2365 445 2399
rect 345 2327 445 2365
rect 503 2399 603 2415
rect 503 2365 519 2399
rect 587 2365 603 2399
rect 503 2327 603 2365
rect 661 2399 761 2415
rect 661 2365 677 2399
rect 745 2365 761 2399
rect 661 2327 761 2365
rect 819 2399 919 2415
rect 819 2365 835 2399
rect 903 2365 919 2399
rect 819 2327 919 2365
rect 977 2399 1077 2415
rect 977 2365 993 2399
rect 1061 2365 1077 2399
rect 977 2327 1077 2365
rect 1135 2399 1235 2415
rect 1135 2365 1151 2399
rect 1219 2365 1235 2399
rect 1135 2327 1235 2365
rect 1293 2399 1393 2415
rect 1293 2365 1309 2399
rect 1377 2365 1393 2399
rect 1293 2327 1393 2365
rect 1451 2399 1551 2415
rect 1451 2365 1467 2399
rect 1535 2365 1551 2399
rect 1451 2327 1551 2365
rect -1551 1289 -1451 1327
rect -1551 1255 -1535 1289
rect -1467 1255 -1451 1289
rect -1551 1239 -1451 1255
rect -1393 1289 -1293 1327
rect -1393 1255 -1377 1289
rect -1309 1255 -1293 1289
rect -1393 1239 -1293 1255
rect -1235 1289 -1135 1327
rect -1235 1255 -1219 1289
rect -1151 1255 -1135 1289
rect -1235 1239 -1135 1255
rect -1077 1289 -977 1327
rect -1077 1255 -1061 1289
rect -993 1255 -977 1289
rect -1077 1239 -977 1255
rect -919 1289 -819 1327
rect -919 1255 -903 1289
rect -835 1255 -819 1289
rect -919 1239 -819 1255
rect -761 1289 -661 1327
rect -761 1255 -745 1289
rect -677 1255 -661 1289
rect -761 1239 -661 1255
rect -603 1289 -503 1327
rect -603 1255 -587 1289
rect -519 1255 -503 1289
rect -603 1239 -503 1255
rect -445 1289 -345 1327
rect -445 1255 -429 1289
rect -361 1255 -345 1289
rect -445 1239 -345 1255
rect -287 1289 -187 1327
rect -287 1255 -271 1289
rect -203 1255 -187 1289
rect -287 1239 -187 1255
rect -129 1289 -29 1327
rect -129 1255 -113 1289
rect -45 1255 -29 1289
rect -129 1239 -29 1255
rect 29 1289 129 1327
rect 29 1255 45 1289
rect 113 1255 129 1289
rect 29 1239 129 1255
rect 187 1289 287 1327
rect 187 1255 203 1289
rect 271 1255 287 1289
rect 187 1239 287 1255
rect 345 1289 445 1327
rect 345 1255 361 1289
rect 429 1255 445 1289
rect 345 1239 445 1255
rect 503 1289 603 1327
rect 503 1255 519 1289
rect 587 1255 603 1289
rect 503 1239 603 1255
rect 661 1289 761 1327
rect 661 1255 677 1289
rect 745 1255 761 1289
rect 661 1239 761 1255
rect 819 1289 919 1327
rect 819 1255 835 1289
rect 903 1255 919 1289
rect 819 1239 919 1255
rect 977 1289 1077 1327
rect 977 1255 993 1289
rect 1061 1255 1077 1289
rect 977 1239 1077 1255
rect 1135 1289 1235 1327
rect 1135 1255 1151 1289
rect 1219 1255 1235 1289
rect 1135 1239 1235 1255
rect 1293 1289 1393 1327
rect 1293 1255 1309 1289
rect 1377 1255 1393 1289
rect 1293 1239 1393 1255
rect 1451 1289 1551 1327
rect 1451 1255 1467 1289
rect 1535 1255 1551 1289
rect 1451 1239 1551 1255
rect -1551 1181 -1451 1197
rect -1551 1147 -1535 1181
rect -1467 1147 -1451 1181
rect -1551 1109 -1451 1147
rect -1393 1181 -1293 1197
rect -1393 1147 -1377 1181
rect -1309 1147 -1293 1181
rect -1393 1109 -1293 1147
rect -1235 1181 -1135 1197
rect -1235 1147 -1219 1181
rect -1151 1147 -1135 1181
rect -1235 1109 -1135 1147
rect -1077 1181 -977 1197
rect -1077 1147 -1061 1181
rect -993 1147 -977 1181
rect -1077 1109 -977 1147
rect -919 1181 -819 1197
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -919 1109 -819 1147
rect -761 1181 -661 1197
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -761 1109 -661 1147
rect -603 1181 -503 1197
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -603 1109 -503 1147
rect -445 1181 -345 1197
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -445 1109 -345 1147
rect -287 1181 -187 1197
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -287 1109 -187 1147
rect -129 1181 -29 1197
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect -129 1109 -29 1147
rect 29 1181 129 1197
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 29 1109 129 1147
rect 187 1181 287 1197
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 187 1109 287 1147
rect 345 1181 445 1197
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 345 1109 445 1147
rect 503 1181 603 1197
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 503 1109 603 1147
rect 661 1181 761 1197
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 661 1109 761 1147
rect 819 1181 919 1197
rect 819 1147 835 1181
rect 903 1147 919 1181
rect 819 1109 919 1147
rect 977 1181 1077 1197
rect 977 1147 993 1181
rect 1061 1147 1077 1181
rect 977 1109 1077 1147
rect 1135 1181 1235 1197
rect 1135 1147 1151 1181
rect 1219 1147 1235 1181
rect 1135 1109 1235 1147
rect 1293 1181 1393 1197
rect 1293 1147 1309 1181
rect 1377 1147 1393 1181
rect 1293 1109 1393 1147
rect 1451 1181 1551 1197
rect 1451 1147 1467 1181
rect 1535 1147 1551 1181
rect 1451 1109 1551 1147
rect -1551 71 -1451 109
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 109
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 109
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 109
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 109
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 109
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 109
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 109
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -109 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -109 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -109 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -109 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -109 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -109 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -109 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -109 1551 -71
rect -1551 -1147 -1451 -1109
rect -1551 -1181 -1535 -1147
rect -1467 -1181 -1451 -1147
rect -1551 -1197 -1451 -1181
rect -1393 -1147 -1293 -1109
rect -1393 -1181 -1377 -1147
rect -1309 -1181 -1293 -1147
rect -1393 -1197 -1293 -1181
rect -1235 -1147 -1135 -1109
rect -1235 -1181 -1219 -1147
rect -1151 -1181 -1135 -1147
rect -1235 -1197 -1135 -1181
rect -1077 -1147 -977 -1109
rect -1077 -1181 -1061 -1147
rect -993 -1181 -977 -1147
rect -1077 -1197 -977 -1181
rect -919 -1147 -819 -1109
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -919 -1197 -819 -1181
rect -761 -1147 -661 -1109
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -761 -1197 -661 -1181
rect -603 -1147 -503 -1109
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -603 -1197 -503 -1181
rect -445 -1147 -345 -1109
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -445 -1197 -345 -1181
rect -287 -1147 -187 -1109
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -287 -1197 -187 -1181
rect -129 -1147 -29 -1109
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect -129 -1197 -29 -1181
rect 29 -1147 129 -1109
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 29 -1197 129 -1181
rect 187 -1147 287 -1109
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 187 -1197 287 -1181
rect 345 -1147 445 -1109
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 345 -1197 445 -1181
rect 503 -1147 603 -1109
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 503 -1197 603 -1181
rect 661 -1147 761 -1109
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 661 -1197 761 -1181
rect 819 -1147 919 -1109
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect 819 -1197 919 -1181
rect 977 -1147 1077 -1109
rect 977 -1181 993 -1147
rect 1061 -1181 1077 -1147
rect 977 -1197 1077 -1181
rect 1135 -1147 1235 -1109
rect 1135 -1181 1151 -1147
rect 1219 -1181 1235 -1147
rect 1135 -1197 1235 -1181
rect 1293 -1147 1393 -1109
rect 1293 -1181 1309 -1147
rect 1377 -1181 1393 -1147
rect 1293 -1197 1393 -1181
rect 1451 -1147 1551 -1109
rect 1451 -1181 1467 -1147
rect 1535 -1181 1551 -1147
rect 1451 -1197 1551 -1181
rect -1551 -1255 -1451 -1239
rect -1551 -1289 -1535 -1255
rect -1467 -1289 -1451 -1255
rect -1551 -1327 -1451 -1289
rect -1393 -1255 -1293 -1239
rect -1393 -1289 -1377 -1255
rect -1309 -1289 -1293 -1255
rect -1393 -1327 -1293 -1289
rect -1235 -1255 -1135 -1239
rect -1235 -1289 -1219 -1255
rect -1151 -1289 -1135 -1255
rect -1235 -1327 -1135 -1289
rect -1077 -1255 -977 -1239
rect -1077 -1289 -1061 -1255
rect -993 -1289 -977 -1255
rect -1077 -1327 -977 -1289
rect -919 -1255 -819 -1239
rect -919 -1289 -903 -1255
rect -835 -1289 -819 -1255
rect -919 -1327 -819 -1289
rect -761 -1255 -661 -1239
rect -761 -1289 -745 -1255
rect -677 -1289 -661 -1255
rect -761 -1327 -661 -1289
rect -603 -1255 -503 -1239
rect -603 -1289 -587 -1255
rect -519 -1289 -503 -1255
rect -603 -1327 -503 -1289
rect -445 -1255 -345 -1239
rect -445 -1289 -429 -1255
rect -361 -1289 -345 -1255
rect -445 -1327 -345 -1289
rect -287 -1255 -187 -1239
rect -287 -1289 -271 -1255
rect -203 -1289 -187 -1255
rect -287 -1327 -187 -1289
rect -129 -1255 -29 -1239
rect -129 -1289 -113 -1255
rect -45 -1289 -29 -1255
rect -129 -1327 -29 -1289
rect 29 -1255 129 -1239
rect 29 -1289 45 -1255
rect 113 -1289 129 -1255
rect 29 -1327 129 -1289
rect 187 -1255 287 -1239
rect 187 -1289 203 -1255
rect 271 -1289 287 -1255
rect 187 -1327 287 -1289
rect 345 -1255 445 -1239
rect 345 -1289 361 -1255
rect 429 -1289 445 -1255
rect 345 -1327 445 -1289
rect 503 -1255 603 -1239
rect 503 -1289 519 -1255
rect 587 -1289 603 -1255
rect 503 -1327 603 -1289
rect 661 -1255 761 -1239
rect 661 -1289 677 -1255
rect 745 -1289 761 -1255
rect 661 -1327 761 -1289
rect 819 -1255 919 -1239
rect 819 -1289 835 -1255
rect 903 -1289 919 -1255
rect 819 -1327 919 -1289
rect 977 -1255 1077 -1239
rect 977 -1289 993 -1255
rect 1061 -1289 1077 -1255
rect 977 -1327 1077 -1289
rect 1135 -1255 1235 -1239
rect 1135 -1289 1151 -1255
rect 1219 -1289 1235 -1255
rect 1135 -1327 1235 -1289
rect 1293 -1255 1393 -1239
rect 1293 -1289 1309 -1255
rect 1377 -1289 1393 -1255
rect 1293 -1327 1393 -1289
rect 1451 -1255 1551 -1239
rect 1451 -1289 1467 -1255
rect 1535 -1289 1551 -1255
rect 1451 -1327 1551 -1289
rect -1551 -2365 -1451 -2327
rect -1551 -2399 -1535 -2365
rect -1467 -2399 -1451 -2365
rect -1551 -2415 -1451 -2399
rect -1393 -2365 -1293 -2327
rect -1393 -2399 -1377 -2365
rect -1309 -2399 -1293 -2365
rect -1393 -2415 -1293 -2399
rect -1235 -2365 -1135 -2327
rect -1235 -2399 -1219 -2365
rect -1151 -2399 -1135 -2365
rect -1235 -2415 -1135 -2399
rect -1077 -2365 -977 -2327
rect -1077 -2399 -1061 -2365
rect -993 -2399 -977 -2365
rect -1077 -2415 -977 -2399
rect -919 -2365 -819 -2327
rect -919 -2399 -903 -2365
rect -835 -2399 -819 -2365
rect -919 -2415 -819 -2399
rect -761 -2365 -661 -2327
rect -761 -2399 -745 -2365
rect -677 -2399 -661 -2365
rect -761 -2415 -661 -2399
rect -603 -2365 -503 -2327
rect -603 -2399 -587 -2365
rect -519 -2399 -503 -2365
rect -603 -2415 -503 -2399
rect -445 -2365 -345 -2327
rect -445 -2399 -429 -2365
rect -361 -2399 -345 -2365
rect -445 -2415 -345 -2399
rect -287 -2365 -187 -2327
rect -287 -2399 -271 -2365
rect -203 -2399 -187 -2365
rect -287 -2415 -187 -2399
rect -129 -2365 -29 -2327
rect -129 -2399 -113 -2365
rect -45 -2399 -29 -2365
rect -129 -2415 -29 -2399
rect 29 -2365 129 -2327
rect 29 -2399 45 -2365
rect 113 -2399 129 -2365
rect 29 -2415 129 -2399
rect 187 -2365 287 -2327
rect 187 -2399 203 -2365
rect 271 -2399 287 -2365
rect 187 -2415 287 -2399
rect 345 -2365 445 -2327
rect 345 -2399 361 -2365
rect 429 -2399 445 -2365
rect 345 -2415 445 -2399
rect 503 -2365 603 -2327
rect 503 -2399 519 -2365
rect 587 -2399 603 -2365
rect 503 -2415 603 -2399
rect 661 -2365 761 -2327
rect 661 -2399 677 -2365
rect 745 -2399 761 -2365
rect 661 -2415 761 -2399
rect 819 -2365 919 -2327
rect 819 -2399 835 -2365
rect 903 -2399 919 -2365
rect 819 -2415 919 -2399
rect 977 -2365 1077 -2327
rect 977 -2399 993 -2365
rect 1061 -2399 1077 -2365
rect 977 -2415 1077 -2399
rect 1135 -2365 1235 -2327
rect 1135 -2399 1151 -2365
rect 1219 -2399 1235 -2365
rect 1135 -2415 1235 -2399
rect 1293 -2365 1393 -2327
rect 1293 -2399 1309 -2365
rect 1377 -2399 1393 -2365
rect 1293 -2415 1393 -2399
rect 1451 -2365 1551 -2327
rect 1451 -2399 1467 -2365
rect 1535 -2399 1551 -2365
rect 1451 -2415 1551 -2399
rect -1551 -2473 -1451 -2457
rect -1551 -2507 -1535 -2473
rect -1467 -2507 -1451 -2473
rect -1551 -2545 -1451 -2507
rect -1393 -2473 -1293 -2457
rect -1393 -2507 -1377 -2473
rect -1309 -2507 -1293 -2473
rect -1393 -2545 -1293 -2507
rect -1235 -2473 -1135 -2457
rect -1235 -2507 -1219 -2473
rect -1151 -2507 -1135 -2473
rect -1235 -2545 -1135 -2507
rect -1077 -2473 -977 -2457
rect -1077 -2507 -1061 -2473
rect -993 -2507 -977 -2473
rect -1077 -2545 -977 -2507
rect -919 -2473 -819 -2457
rect -919 -2507 -903 -2473
rect -835 -2507 -819 -2473
rect -919 -2545 -819 -2507
rect -761 -2473 -661 -2457
rect -761 -2507 -745 -2473
rect -677 -2507 -661 -2473
rect -761 -2545 -661 -2507
rect -603 -2473 -503 -2457
rect -603 -2507 -587 -2473
rect -519 -2507 -503 -2473
rect -603 -2545 -503 -2507
rect -445 -2473 -345 -2457
rect -445 -2507 -429 -2473
rect -361 -2507 -345 -2473
rect -445 -2545 -345 -2507
rect -287 -2473 -187 -2457
rect -287 -2507 -271 -2473
rect -203 -2507 -187 -2473
rect -287 -2545 -187 -2507
rect -129 -2473 -29 -2457
rect -129 -2507 -113 -2473
rect -45 -2507 -29 -2473
rect -129 -2545 -29 -2507
rect 29 -2473 129 -2457
rect 29 -2507 45 -2473
rect 113 -2507 129 -2473
rect 29 -2545 129 -2507
rect 187 -2473 287 -2457
rect 187 -2507 203 -2473
rect 271 -2507 287 -2473
rect 187 -2545 287 -2507
rect 345 -2473 445 -2457
rect 345 -2507 361 -2473
rect 429 -2507 445 -2473
rect 345 -2545 445 -2507
rect 503 -2473 603 -2457
rect 503 -2507 519 -2473
rect 587 -2507 603 -2473
rect 503 -2545 603 -2507
rect 661 -2473 761 -2457
rect 661 -2507 677 -2473
rect 745 -2507 761 -2473
rect 661 -2545 761 -2507
rect 819 -2473 919 -2457
rect 819 -2507 835 -2473
rect 903 -2507 919 -2473
rect 819 -2545 919 -2507
rect 977 -2473 1077 -2457
rect 977 -2507 993 -2473
rect 1061 -2507 1077 -2473
rect 977 -2545 1077 -2507
rect 1135 -2473 1235 -2457
rect 1135 -2507 1151 -2473
rect 1219 -2507 1235 -2473
rect 1135 -2545 1235 -2507
rect 1293 -2473 1393 -2457
rect 1293 -2507 1309 -2473
rect 1377 -2507 1393 -2473
rect 1293 -2545 1393 -2507
rect 1451 -2473 1551 -2457
rect 1451 -2507 1467 -2473
rect 1535 -2507 1551 -2473
rect 1451 -2545 1551 -2507
rect -1551 -3583 -1451 -3545
rect -1551 -3617 -1535 -3583
rect -1467 -3617 -1451 -3583
rect -1551 -3633 -1451 -3617
rect -1393 -3583 -1293 -3545
rect -1393 -3617 -1377 -3583
rect -1309 -3617 -1293 -3583
rect -1393 -3633 -1293 -3617
rect -1235 -3583 -1135 -3545
rect -1235 -3617 -1219 -3583
rect -1151 -3617 -1135 -3583
rect -1235 -3633 -1135 -3617
rect -1077 -3583 -977 -3545
rect -1077 -3617 -1061 -3583
rect -993 -3617 -977 -3583
rect -1077 -3633 -977 -3617
rect -919 -3583 -819 -3545
rect -919 -3617 -903 -3583
rect -835 -3617 -819 -3583
rect -919 -3633 -819 -3617
rect -761 -3583 -661 -3545
rect -761 -3617 -745 -3583
rect -677 -3617 -661 -3583
rect -761 -3633 -661 -3617
rect -603 -3583 -503 -3545
rect -603 -3617 -587 -3583
rect -519 -3617 -503 -3583
rect -603 -3633 -503 -3617
rect -445 -3583 -345 -3545
rect -445 -3617 -429 -3583
rect -361 -3617 -345 -3583
rect -445 -3633 -345 -3617
rect -287 -3583 -187 -3545
rect -287 -3617 -271 -3583
rect -203 -3617 -187 -3583
rect -287 -3633 -187 -3617
rect -129 -3583 -29 -3545
rect -129 -3617 -113 -3583
rect -45 -3617 -29 -3583
rect -129 -3633 -29 -3617
rect 29 -3583 129 -3545
rect 29 -3617 45 -3583
rect 113 -3617 129 -3583
rect 29 -3633 129 -3617
rect 187 -3583 287 -3545
rect 187 -3617 203 -3583
rect 271 -3617 287 -3583
rect 187 -3633 287 -3617
rect 345 -3583 445 -3545
rect 345 -3617 361 -3583
rect 429 -3617 445 -3583
rect 345 -3633 445 -3617
rect 503 -3583 603 -3545
rect 503 -3617 519 -3583
rect 587 -3617 603 -3583
rect 503 -3633 603 -3617
rect 661 -3583 761 -3545
rect 661 -3617 677 -3583
rect 745 -3617 761 -3583
rect 661 -3633 761 -3617
rect 819 -3583 919 -3545
rect 819 -3617 835 -3583
rect 903 -3617 919 -3583
rect 819 -3633 919 -3617
rect 977 -3583 1077 -3545
rect 977 -3617 993 -3583
rect 1061 -3617 1077 -3583
rect 977 -3633 1077 -3617
rect 1135 -3583 1235 -3545
rect 1135 -3617 1151 -3583
rect 1219 -3617 1235 -3583
rect 1135 -3633 1235 -3617
rect 1293 -3583 1393 -3545
rect 1293 -3617 1309 -3583
rect 1377 -3617 1393 -3583
rect 1293 -3633 1393 -3617
rect 1451 -3583 1551 -3545
rect 1451 -3617 1467 -3583
rect 1535 -3617 1551 -3583
rect 1451 -3633 1551 -3617
rect -1551 -3691 -1451 -3675
rect -1551 -3725 -1535 -3691
rect -1467 -3725 -1451 -3691
rect -1551 -3763 -1451 -3725
rect -1393 -3691 -1293 -3675
rect -1393 -3725 -1377 -3691
rect -1309 -3725 -1293 -3691
rect -1393 -3763 -1293 -3725
rect -1235 -3691 -1135 -3675
rect -1235 -3725 -1219 -3691
rect -1151 -3725 -1135 -3691
rect -1235 -3763 -1135 -3725
rect -1077 -3691 -977 -3675
rect -1077 -3725 -1061 -3691
rect -993 -3725 -977 -3691
rect -1077 -3763 -977 -3725
rect -919 -3691 -819 -3675
rect -919 -3725 -903 -3691
rect -835 -3725 -819 -3691
rect -919 -3763 -819 -3725
rect -761 -3691 -661 -3675
rect -761 -3725 -745 -3691
rect -677 -3725 -661 -3691
rect -761 -3763 -661 -3725
rect -603 -3691 -503 -3675
rect -603 -3725 -587 -3691
rect -519 -3725 -503 -3691
rect -603 -3763 -503 -3725
rect -445 -3691 -345 -3675
rect -445 -3725 -429 -3691
rect -361 -3725 -345 -3691
rect -445 -3763 -345 -3725
rect -287 -3691 -187 -3675
rect -287 -3725 -271 -3691
rect -203 -3725 -187 -3691
rect -287 -3763 -187 -3725
rect -129 -3691 -29 -3675
rect -129 -3725 -113 -3691
rect -45 -3725 -29 -3691
rect -129 -3763 -29 -3725
rect 29 -3691 129 -3675
rect 29 -3725 45 -3691
rect 113 -3725 129 -3691
rect 29 -3763 129 -3725
rect 187 -3691 287 -3675
rect 187 -3725 203 -3691
rect 271 -3725 287 -3691
rect 187 -3763 287 -3725
rect 345 -3691 445 -3675
rect 345 -3725 361 -3691
rect 429 -3725 445 -3691
rect 345 -3763 445 -3725
rect 503 -3691 603 -3675
rect 503 -3725 519 -3691
rect 587 -3725 603 -3691
rect 503 -3763 603 -3725
rect 661 -3691 761 -3675
rect 661 -3725 677 -3691
rect 745 -3725 761 -3691
rect 661 -3763 761 -3725
rect 819 -3691 919 -3675
rect 819 -3725 835 -3691
rect 903 -3725 919 -3691
rect 819 -3763 919 -3725
rect 977 -3691 1077 -3675
rect 977 -3725 993 -3691
rect 1061 -3725 1077 -3691
rect 977 -3763 1077 -3725
rect 1135 -3691 1235 -3675
rect 1135 -3725 1151 -3691
rect 1219 -3725 1235 -3691
rect 1135 -3763 1235 -3725
rect 1293 -3691 1393 -3675
rect 1293 -3725 1309 -3691
rect 1377 -3725 1393 -3691
rect 1293 -3763 1393 -3725
rect 1451 -3691 1551 -3675
rect 1451 -3725 1467 -3691
rect 1535 -3725 1551 -3691
rect 1451 -3763 1551 -3725
rect -1551 -4801 -1451 -4763
rect -1551 -4835 -1535 -4801
rect -1467 -4835 -1451 -4801
rect -1551 -4851 -1451 -4835
rect -1393 -4801 -1293 -4763
rect -1393 -4835 -1377 -4801
rect -1309 -4835 -1293 -4801
rect -1393 -4851 -1293 -4835
rect -1235 -4801 -1135 -4763
rect -1235 -4835 -1219 -4801
rect -1151 -4835 -1135 -4801
rect -1235 -4851 -1135 -4835
rect -1077 -4801 -977 -4763
rect -1077 -4835 -1061 -4801
rect -993 -4835 -977 -4801
rect -1077 -4851 -977 -4835
rect -919 -4801 -819 -4763
rect -919 -4835 -903 -4801
rect -835 -4835 -819 -4801
rect -919 -4851 -819 -4835
rect -761 -4801 -661 -4763
rect -761 -4835 -745 -4801
rect -677 -4835 -661 -4801
rect -761 -4851 -661 -4835
rect -603 -4801 -503 -4763
rect -603 -4835 -587 -4801
rect -519 -4835 -503 -4801
rect -603 -4851 -503 -4835
rect -445 -4801 -345 -4763
rect -445 -4835 -429 -4801
rect -361 -4835 -345 -4801
rect -445 -4851 -345 -4835
rect -287 -4801 -187 -4763
rect -287 -4835 -271 -4801
rect -203 -4835 -187 -4801
rect -287 -4851 -187 -4835
rect -129 -4801 -29 -4763
rect -129 -4835 -113 -4801
rect -45 -4835 -29 -4801
rect -129 -4851 -29 -4835
rect 29 -4801 129 -4763
rect 29 -4835 45 -4801
rect 113 -4835 129 -4801
rect 29 -4851 129 -4835
rect 187 -4801 287 -4763
rect 187 -4835 203 -4801
rect 271 -4835 287 -4801
rect 187 -4851 287 -4835
rect 345 -4801 445 -4763
rect 345 -4835 361 -4801
rect 429 -4835 445 -4801
rect 345 -4851 445 -4835
rect 503 -4801 603 -4763
rect 503 -4835 519 -4801
rect 587 -4835 603 -4801
rect 503 -4851 603 -4835
rect 661 -4801 761 -4763
rect 661 -4835 677 -4801
rect 745 -4835 761 -4801
rect 661 -4851 761 -4835
rect 819 -4801 919 -4763
rect 819 -4835 835 -4801
rect 903 -4835 919 -4801
rect 819 -4851 919 -4835
rect 977 -4801 1077 -4763
rect 977 -4835 993 -4801
rect 1061 -4835 1077 -4801
rect 977 -4851 1077 -4835
rect 1135 -4801 1235 -4763
rect 1135 -4835 1151 -4801
rect 1219 -4835 1235 -4801
rect 1135 -4851 1235 -4835
rect 1293 -4801 1393 -4763
rect 1293 -4835 1309 -4801
rect 1377 -4835 1393 -4801
rect 1293 -4851 1393 -4835
rect 1451 -4801 1551 -4763
rect 1451 -4835 1467 -4801
rect 1535 -4835 1551 -4801
rect 1451 -4851 1551 -4835
rect -1551 -4909 -1451 -4893
rect -1551 -4943 -1535 -4909
rect -1467 -4943 -1451 -4909
rect -1551 -4981 -1451 -4943
rect -1393 -4909 -1293 -4893
rect -1393 -4943 -1377 -4909
rect -1309 -4943 -1293 -4909
rect -1393 -4981 -1293 -4943
rect -1235 -4909 -1135 -4893
rect -1235 -4943 -1219 -4909
rect -1151 -4943 -1135 -4909
rect -1235 -4981 -1135 -4943
rect -1077 -4909 -977 -4893
rect -1077 -4943 -1061 -4909
rect -993 -4943 -977 -4909
rect -1077 -4981 -977 -4943
rect -919 -4909 -819 -4893
rect -919 -4943 -903 -4909
rect -835 -4943 -819 -4909
rect -919 -4981 -819 -4943
rect -761 -4909 -661 -4893
rect -761 -4943 -745 -4909
rect -677 -4943 -661 -4909
rect -761 -4981 -661 -4943
rect -603 -4909 -503 -4893
rect -603 -4943 -587 -4909
rect -519 -4943 -503 -4909
rect -603 -4981 -503 -4943
rect -445 -4909 -345 -4893
rect -445 -4943 -429 -4909
rect -361 -4943 -345 -4909
rect -445 -4981 -345 -4943
rect -287 -4909 -187 -4893
rect -287 -4943 -271 -4909
rect -203 -4943 -187 -4909
rect -287 -4981 -187 -4943
rect -129 -4909 -29 -4893
rect -129 -4943 -113 -4909
rect -45 -4943 -29 -4909
rect -129 -4981 -29 -4943
rect 29 -4909 129 -4893
rect 29 -4943 45 -4909
rect 113 -4943 129 -4909
rect 29 -4981 129 -4943
rect 187 -4909 287 -4893
rect 187 -4943 203 -4909
rect 271 -4943 287 -4909
rect 187 -4981 287 -4943
rect 345 -4909 445 -4893
rect 345 -4943 361 -4909
rect 429 -4943 445 -4909
rect 345 -4981 445 -4943
rect 503 -4909 603 -4893
rect 503 -4943 519 -4909
rect 587 -4943 603 -4909
rect 503 -4981 603 -4943
rect 661 -4909 761 -4893
rect 661 -4943 677 -4909
rect 745 -4943 761 -4909
rect 661 -4981 761 -4943
rect 819 -4909 919 -4893
rect 819 -4943 835 -4909
rect 903 -4943 919 -4909
rect 819 -4981 919 -4943
rect 977 -4909 1077 -4893
rect 977 -4943 993 -4909
rect 1061 -4943 1077 -4909
rect 977 -4981 1077 -4943
rect 1135 -4909 1235 -4893
rect 1135 -4943 1151 -4909
rect 1219 -4943 1235 -4909
rect 1135 -4981 1235 -4943
rect 1293 -4909 1393 -4893
rect 1293 -4943 1309 -4909
rect 1377 -4943 1393 -4909
rect 1293 -4981 1393 -4943
rect 1451 -4909 1551 -4893
rect 1451 -4943 1467 -4909
rect 1535 -4943 1551 -4909
rect 1451 -4981 1551 -4943
rect -1551 -6019 -1451 -5981
rect -1551 -6053 -1535 -6019
rect -1467 -6053 -1451 -6019
rect -1551 -6069 -1451 -6053
rect -1393 -6019 -1293 -5981
rect -1393 -6053 -1377 -6019
rect -1309 -6053 -1293 -6019
rect -1393 -6069 -1293 -6053
rect -1235 -6019 -1135 -5981
rect -1235 -6053 -1219 -6019
rect -1151 -6053 -1135 -6019
rect -1235 -6069 -1135 -6053
rect -1077 -6019 -977 -5981
rect -1077 -6053 -1061 -6019
rect -993 -6053 -977 -6019
rect -1077 -6069 -977 -6053
rect -919 -6019 -819 -5981
rect -919 -6053 -903 -6019
rect -835 -6053 -819 -6019
rect -919 -6069 -819 -6053
rect -761 -6019 -661 -5981
rect -761 -6053 -745 -6019
rect -677 -6053 -661 -6019
rect -761 -6069 -661 -6053
rect -603 -6019 -503 -5981
rect -603 -6053 -587 -6019
rect -519 -6053 -503 -6019
rect -603 -6069 -503 -6053
rect -445 -6019 -345 -5981
rect -445 -6053 -429 -6019
rect -361 -6053 -345 -6019
rect -445 -6069 -345 -6053
rect -287 -6019 -187 -5981
rect -287 -6053 -271 -6019
rect -203 -6053 -187 -6019
rect -287 -6069 -187 -6053
rect -129 -6019 -29 -5981
rect -129 -6053 -113 -6019
rect -45 -6053 -29 -6019
rect -129 -6069 -29 -6053
rect 29 -6019 129 -5981
rect 29 -6053 45 -6019
rect 113 -6053 129 -6019
rect 29 -6069 129 -6053
rect 187 -6019 287 -5981
rect 187 -6053 203 -6019
rect 271 -6053 287 -6019
rect 187 -6069 287 -6053
rect 345 -6019 445 -5981
rect 345 -6053 361 -6019
rect 429 -6053 445 -6019
rect 345 -6069 445 -6053
rect 503 -6019 603 -5981
rect 503 -6053 519 -6019
rect 587 -6053 603 -6019
rect 503 -6069 603 -6053
rect 661 -6019 761 -5981
rect 661 -6053 677 -6019
rect 745 -6053 761 -6019
rect 661 -6069 761 -6053
rect 819 -6019 919 -5981
rect 819 -6053 835 -6019
rect 903 -6053 919 -6019
rect 819 -6069 919 -6053
rect 977 -6019 1077 -5981
rect 977 -6053 993 -6019
rect 1061 -6053 1077 -6019
rect 977 -6069 1077 -6053
rect 1135 -6019 1235 -5981
rect 1135 -6053 1151 -6019
rect 1219 -6053 1235 -6019
rect 1135 -6069 1235 -6053
rect 1293 -6019 1393 -5981
rect 1293 -6053 1309 -6019
rect 1377 -6053 1393 -6019
rect 1293 -6069 1393 -6053
rect 1451 -6019 1551 -5981
rect 1451 -6053 1467 -6019
rect 1535 -6053 1551 -6019
rect 1451 -6069 1551 -6053
<< polycont >>
rect -1535 6019 -1467 6053
rect -1377 6019 -1309 6053
rect -1219 6019 -1151 6053
rect -1061 6019 -993 6053
rect -903 6019 -835 6053
rect -745 6019 -677 6053
rect -587 6019 -519 6053
rect -429 6019 -361 6053
rect -271 6019 -203 6053
rect -113 6019 -45 6053
rect 45 6019 113 6053
rect 203 6019 271 6053
rect 361 6019 429 6053
rect 519 6019 587 6053
rect 677 6019 745 6053
rect 835 6019 903 6053
rect 993 6019 1061 6053
rect 1151 6019 1219 6053
rect 1309 6019 1377 6053
rect 1467 6019 1535 6053
rect -1535 4909 -1467 4943
rect -1377 4909 -1309 4943
rect -1219 4909 -1151 4943
rect -1061 4909 -993 4943
rect -903 4909 -835 4943
rect -745 4909 -677 4943
rect -587 4909 -519 4943
rect -429 4909 -361 4943
rect -271 4909 -203 4943
rect -113 4909 -45 4943
rect 45 4909 113 4943
rect 203 4909 271 4943
rect 361 4909 429 4943
rect 519 4909 587 4943
rect 677 4909 745 4943
rect 835 4909 903 4943
rect 993 4909 1061 4943
rect 1151 4909 1219 4943
rect 1309 4909 1377 4943
rect 1467 4909 1535 4943
rect -1535 4801 -1467 4835
rect -1377 4801 -1309 4835
rect -1219 4801 -1151 4835
rect -1061 4801 -993 4835
rect -903 4801 -835 4835
rect -745 4801 -677 4835
rect -587 4801 -519 4835
rect -429 4801 -361 4835
rect -271 4801 -203 4835
rect -113 4801 -45 4835
rect 45 4801 113 4835
rect 203 4801 271 4835
rect 361 4801 429 4835
rect 519 4801 587 4835
rect 677 4801 745 4835
rect 835 4801 903 4835
rect 993 4801 1061 4835
rect 1151 4801 1219 4835
rect 1309 4801 1377 4835
rect 1467 4801 1535 4835
rect -1535 3691 -1467 3725
rect -1377 3691 -1309 3725
rect -1219 3691 -1151 3725
rect -1061 3691 -993 3725
rect -903 3691 -835 3725
rect -745 3691 -677 3725
rect -587 3691 -519 3725
rect -429 3691 -361 3725
rect -271 3691 -203 3725
rect -113 3691 -45 3725
rect 45 3691 113 3725
rect 203 3691 271 3725
rect 361 3691 429 3725
rect 519 3691 587 3725
rect 677 3691 745 3725
rect 835 3691 903 3725
rect 993 3691 1061 3725
rect 1151 3691 1219 3725
rect 1309 3691 1377 3725
rect 1467 3691 1535 3725
rect -1535 3583 -1467 3617
rect -1377 3583 -1309 3617
rect -1219 3583 -1151 3617
rect -1061 3583 -993 3617
rect -903 3583 -835 3617
rect -745 3583 -677 3617
rect -587 3583 -519 3617
rect -429 3583 -361 3617
rect -271 3583 -203 3617
rect -113 3583 -45 3617
rect 45 3583 113 3617
rect 203 3583 271 3617
rect 361 3583 429 3617
rect 519 3583 587 3617
rect 677 3583 745 3617
rect 835 3583 903 3617
rect 993 3583 1061 3617
rect 1151 3583 1219 3617
rect 1309 3583 1377 3617
rect 1467 3583 1535 3617
rect -1535 2473 -1467 2507
rect -1377 2473 -1309 2507
rect -1219 2473 -1151 2507
rect -1061 2473 -993 2507
rect -903 2473 -835 2507
rect -745 2473 -677 2507
rect -587 2473 -519 2507
rect -429 2473 -361 2507
rect -271 2473 -203 2507
rect -113 2473 -45 2507
rect 45 2473 113 2507
rect 203 2473 271 2507
rect 361 2473 429 2507
rect 519 2473 587 2507
rect 677 2473 745 2507
rect 835 2473 903 2507
rect 993 2473 1061 2507
rect 1151 2473 1219 2507
rect 1309 2473 1377 2507
rect 1467 2473 1535 2507
rect -1535 2365 -1467 2399
rect -1377 2365 -1309 2399
rect -1219 2365 -1151 2399
rect -1061 2365 -993 2399
rect -903 2365 -835 2399
rect -745 2365 -677 2399
rect -587 2365 -519 2399
rect -429 2365 -361 2399
rect -271 2365 -203 2399
rect -113 2365 -45 2399
rect 45 2365 113 2399
rect 203 2365 271 2399
rect 361 2365 429 2399
rect 519 2365 587 2399
rect 677 2365 745 2399
rect 835 2365 903 2399
rect 993 2365 1061 2399
rect 1151 2365 1219 2399
rect 1309 2365 1377 2399
rect 1467 2365 1535 2399
rect -1535 1255 -1467 1289
rect -1377 1255 -1309 1289
rect -1219 1255 -1151 1289
rect -1061 1255 -993 1289
rect -903 1255 -835 1289
rect -745 1255 -677 1289
rect -587 1255 -519 1289
rect -429 1255 -361 1289
rect -271 1255 -203 1289
rect -113 1255 -45 1289
rect 45 1255 113 1289
rect 203 1255 271 1289
rect 361 1255 429 1289
rect 519 1255 587 1289
rect 677 1255 745 1289
rect 835 1255 903 1289
rect 993 1255 1061 1289
rect 1151 1255 1219 1289
rect 1309 1255 1377 1289
rect 1467 1255 1535 1289
rect -1535 1147 -1467 1181
rect -1377 1147 -1309 1181
rect -1219 1147 -1151 1181
rect -1061 1147 -993 1181
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect 993 1147 1061 1181
rect 1151 1147 1219 1181
rect 1309 1147 1377 1181
rect 1467 1147 1535 1181
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect -1535 -1181 -1467 -1147
rect -1377 -1181 -1309 -1147
rect -1219 -1181 -1151 -1147
rect -1061 -1181 -993 -1147
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
rect 993 -1181 1061 -1147
rect 1151 -1181 1219 -1147
rect 1309 -1181 1377 -1147
rect 1467 -1181 1535 -1147
rect -1535 -1289 -1467 -1255
rect -1377 -1289 -1309 -1255
rect -1219 -1289 -1151 -1255
rect -1061 -1289 -993 -1255
rect -903 -1289 -835 -1255
rect -745 -1289 -677 -1255
rect -587 -1289 -519 -1255
rect -429 -1289 -361 -1255
rect -271 -1289 -203 -1255
rect -113 -1289 -45 -1255
rect 45 -1289 113 -1255
rect 203 -1289 271 -1255
rect 361 -1289 429 -1255
rect 519 -1289 587 -1255
rect 677 -1289 745 -1255
rect 835 -1289 903 -1255
rect 993 -1289 1061 -1255
rect 1151 -1289 1219 -1255
rect 1309 -1289 1377 -1255
rect 1467 -1289 1535 -1255
rect -1535 -2399 -1467 -2365
rect -1377 -2399 -1309 -2365
rect -1219 -2399 -1151 -2365
rect -1061 -2399 -993 -2365
rect -903 -2399 -835 -2365
rect -745 -2399 -677 -2365
rect -587 -2399 -519 -2365
rect -429 -2399 -361 -2365
rect -271 -2399 -203 -2365
rect -113 -2399 -45 -2365
rect 45 -2399 113 -2365
rect 203 -2399 271 -2365
rect 361 -2399 429 -2365
rect 519 -2399 587 -2365
rect 677 -2399 745 -2365
rect 835 -2399 903 -2365
rect 993 -2399 1061 -2365
rect 1151 -2399 1219 -2365
rect 1309 -2399 1377 -2365
rect 1467 -2399 1535 -2365
rect -1535 -2507 -1467 -2473
rect -1377 -2507 -1309 -2473
rect -1219 -2507 -1151 -2473
rect -1061 -2507 -993 -2473
rect -903 -2507 -835 -2473
rect -745 -2507 -677 -2473
rect -587 -2507 -519 -2473
rect -429 -2507 -361 -2473
rect -271 -2507 -203 -2473
rect -113 -2507 -45 -2473
rect 45 -2507 113 -2473
rect 203 -2507 271 -2473
rect 361 -2507 429 -2473
rect 519 -2507 587 -2473
rect 677 -2507 745 -2473
rect 835 -2507 903 -2473
rect 993 -2507 1061 -2473
rect 1151 -2507 1219 -2473
rect 1309 -2507 1377 -2473
rect 1467 -2507 1535 -2473
rect -1535 -3617 -1467 -3583
rect -1377 -3617 -1309 -3583
rect -1219 -3617 -1151 -3583
rect -1061 -3617 -993 -3583
rect -903 -3617 -835 -3583
rect -745 -3617 -677 -3583
rect -587 -3617 -519 -3583
rect -429 -3617 -361 -3583
rect -271 -3617 -203 -3583
rect -113 -3617 -45 -3583
rect 45 -3617 113 -3583
rect 203 -3617 271 -3583
rect 361 -3617 429 -3583
rect 519 -3617 587 -3583
rect 677 -3617 745 -3583
rect 835 -3617 903 -3583
rect 993 -3617 1061 -3583
rect 1151 -3617 1219 -3583
rect 1309 -3617 1377 -3583
rect 1467 -3617 1535 -3583
rect -1535 -3725 -1467 -3691
rect -1377 -3725 -1309 -3691
rect -1219 -3725 -1151 -3691
rect -1061 -3725 -993 -3691
rect -903 -3725 -835 -3691
rect -745 -3725 -677 -3691
rect -587 -3725 -519 -3691
rect -429 -3725 -361 -3691
rect -271 -3725 -203 -3691
rect -113 -3725 -45 -3691
rect 45 -3725 113 -3691
rect 203 -3725 271 -3691
rect 361 -3725 429 -3691
rect 519 -3725 587 -3691
rect 677 -3725 745 -3691
rect 835 -3725 903 -3691
rect 993 -3725 1061 -3691
rect 1151 -3725 1219 -3691
rect 1309 -3725 1377 -3691
rect 1467 -3725 1535 -3691
rect -1535 -4835 -1467 -4801
rect -1377 -4835 -1309 -4801
rect -1219 -4835 -1151 -4801
rect -1061 -4835 -993 -4801
rect -903 -4835 -835 -4801
rect -745 -4835 -677 -4801
rect -587 -4835 -519 -4801
rect -429 -4835 -361 -4801
rect -271 -4835 -203 -4801
rect -113 -4835 -45 -4801
rect 45 -4835 113 -4801
rect 203 -4835 271 -4801
rect 361 -4835 429 -4801
rect 519 -4835 587 -4801
rect 677 -4835 745 -4801
rect 835 -4835 903 -4801
rect 993 -4835 1061 -4801
rect 1151 -4835 1219 -4801
rect 1309 -4835 1377 -4801
rect 1467 -4835 1535 -4801
rect -1535 -4943 -1467 -4909
rect -1377 -4943 -1309 -4909
rect -1219 -4943 -1151 -4909
rect -1061 -4943 -993 -4909
rect -903 -4943 -835 -4909
rect -745 -4943 -677 -4909
rect -587 -4943 -519 -4909
rect -429 -4943 -361 -4909
rect -271 -4943 -203 -4909
rect -113 -4943 -45 -4909
rect 45 -4943 113 -4909
rect 203 -4943 271 -4909
rect 361 -4943 429 -4909
rect 519 -4943 587 -4909
rect 677 -4943 745 -4909
rect 835 -4943 903 -4909
rect 993 -4943 1061 -4909
rect 1151 -4943 1219 -4909
rect 1309 -4943 1377 -4909
rect 1467 -4943 1535 -4909
rect -1535 -6053 -1467 -6019
rect -1377 -6053 -1309 -6019
rect -1219 -6053 -1151 -6019
rect -1061 -6053 -993 -6019
rect -903 -6053 -835 -6019
rect -745 -6053 -677 -6019
rect -587 -6053 -519 -6019
rect -429 -6053 -361 -6019
rect -271 -6053 -203 -6019
rect -113 -6053 -45 -6019
rect 45 -6053 113 -6019
rect 203 -6053 271 -6019
rect 361 -6053 429 -6019
rect 519 -6053 587 -6019
rect 677 -6053 745 -6019
rect 835 -6053 903 -6019
rect 993 -6053 1061 -6019
rect 1151 -6053 1219 -6019
rect 1309 -6053 1377 -6019
rect 1467 -6053 1535 -6019
<< locali >>
rect -1741 6157 -1645 6191
rect 1645 6157 1741 6191
rect -1741 6095 -1707 6157
rect 1707 6095 1741 6157
rect -1551 6019 -1535 6053
rect -1467 6019 -1451 6053
rect -1393 6019 -1377 6053
rect -1309 6019 -1293 6053
rect -1235 6019 -1219 6053
rect -1151 6019 -1135 6053
rect -1077 6019 -1061 6053
rect -993 6019 -977 6053
rect -919 6019 -903 6053
rect -835 6019 -819 6053
rect -761 6019 -745 6053
rect -677 6019 -661 6053
rect -603 6019 -587 6053
rect -519 6019 -503 6053
rect -445 6019 -429 6053
rect -361 6019 -345 6053
rect -287 6019 -271 6053
rect -203 6019 -187 6053
rect -129 6019 -113 6053
rect -45 6019 -29 6053
rect 29 6019 45 6053
rect 113 6019 129 6053
rect 187 6019 203 6053
rect 271 6019 287 6053
rect 345 6019 361 6053
rect 429 6019 445 6053
rect 503 6019 519 6053
rect 587 6019 603 6053
rect 661 6019 677 6053
rect 745 6019 761 6053
rect 819 6019 835 6053
rect 903 6019 919 6053
rect 977 6019 993 6053
rect 1061 6019 1077 6053
rect 1135 6019 1151 6053
rect 1219 6019 1235 6053
rect 1293 6019 1309 6053
rect 1377 6019 1393 6053
rect 1451 6019 1467 6053
rect 1535 6019 1551 6053
rect -1597 5969 -1563 5985
rect -1597 4977 -1563 4993
rect -1439 5969 -1405 5985
rect -1439 4977 -1405 4993
rect -1281 5969 -1247 5985
rect -1281 4977 -1247 4993
rect -1123 5969 -1089 5985
rect -1123 4977 -1089 4993
rect -965 5969 -931 5985
rect -965 4977 -931 4993
rect -807 5969 -773 5985
rect -807 4977 -773 4993
rect -649 5969 -615 5985
rect -649 4977 -615 4993
rect -491 5969 -457 5985
rect -491 4977 -457 4993
rect -333 5969 -299 5985
rect -333 4977 -299 4993
rect -175 5969 -141 5985
rect -175 4977 -141 4993
rect -17 5969 17 5985
rect -17 4977 17 4993
rect 141 5969 175 5985
rect 141 4977 175 4993
rect 299 5969 333 5985
rect 299 4977 333 4993
rect 457 5969 491 5985
rect 457 4977 491 4993
rect 615 5969 649 5985
rect 615 4977 649 4993
rect 773 5969 807 5985
rect 773 4977 807 4993
rect 931 5969 965 5985
rect 931 4977 965 4993
rect 1089 5969 1123 5985
rect 1089 4977 1123 4993
rect 1247 5969 1281 5985
rect 1247 4977 1281 4993
rect 1405 5969 1439 5985
rect 1405 4977 1439 4993
rect 1563 5969 1597 5985
rect 1563 4977 1597 4993
rect -1551 4909 -1535 4943
rect -1467 4909 -1451 4943
rect -1393 4909 -1377 4943
rect -1309 4909 -1293 4943
rect -1235 4909 -1219 4943
rect -1151 4909 -1135 4943
rect -1077 4909 -1061 4943
rect -993 4909 -977 4943
rect -919 4909 -903 4943
rect -835 4909 -819 4943
rect -761 4909 -745 4943
rect -677 4909 -661 4943
rect -603 4909 -587 4943
rect -519 4909 -503 4943
rect -445 4909 -429 4943
rect -361 4909 -345 4943
rect -287 4909 -271 4943
rect -203 4909 -187 4943
rect -129 4909 -113 4943
rect -45 4909 -29 4943
rect 29 4909 45 4943
rect 113 4909 129 4943
rect 187 4909 203 4943
rect 271 4909 287 4943
rect 345 4909 361 4943
rect 429 4909 445 4943
rect 503 4909 519 4943
rect 587 4909 603 4943
rect 661 4909 677 4943
rect 745 4909 761 4943
rect 819 4909 835 4943
rect 903 4909 919 4943
rect 977 4909 993 4943
rect 1061 4909 1077 4943
rect 1135 4909 1151 4943
rect 1219 4909 1235 4943
rect 1293 4909 1309 4943
rect 1377 4909 1393 4943
rect 1451 4909 1467 4943
rect 1535 4909 1551 4943
rect -1551 4801 -1535 4835
rect -1467 4801 -1451 4835
rect -1393 4801 -1377 4835
rect -1309 4801 -1293 4835
rect -1235 4801 -1219 4835
rect -1151 4801 -1135 4835
rect -1077 4801 -1061 4835
rect -993 4801 -977 4835
rect -919 4801 -903 4835
rect -835 4801 -819 4835
rect -761 4801 -745 4835
rect -677 4801 -661 4835
rect -603 4801 -587 4835
rect -519 4801 -503 4835
rect -445 4801 -429 4835
rect -361 4801 -345 4835
rect -287 4801 -271 4835
rect -203 4801 -187 4835
rect -129 4801 -113 4835
rect -45 4801 -29 4835
rect 29 4801 45 4835
rect 113 4801 129 4835
rect 187 4801 203 4835
rect 271 4801 287 4835
rect 345 4801 361 4835
rect 429 4801 445 4835
rect 503 4801 519 4835
rect 587 4801 603 4835
rect 661 4801 677 4835
rect 745 4801 761 4835
rect 819 4801 835 4835
rect 903 4801 919 4835
rect 977 4801 993 4835
rect 1061 4801 1077 4835
rect 1135 4801 1151 4835
rect 1219 4801 1235 4835
rect 1293 4801 1309 4835
rect 1377 4801 1393 4835
rect 1451 4801 1467 4835
rect 1535 4801 1551 4835
rect -1597 4751 -1563 4767
rect -1597 3759 -1563 3775
rect -1439 4751 -1405 4767
rect -1439 3759 -1405 3775
rect -1281 4751 -1247 4767
rect -1281 3759 -1247 3775
rect -1123 4751 -1089 4767
rect -1123 3759 -1089 3775
rect -965 4751 -931 4767
rect -965 3759 -931 3775
rect -807 4751 -773 4767
rect -807 3759 -773 3775
rect -649 4751 -615 4767
rect -649 3759 -615 3775
rect -491 4751 -457 4767
rect -491 3759 -457 3775
rect -333 4751 -299 4767
rect -333 3759 -299 3775
rect -175 4751 -141 4767
rect -175 3759 -141 3775
rect -17 4751 17 4767
rect -17 3759 17 3775
rect 141 4751 175 4767
rect 141 3759 175 3775
rect 299 4751 333 4767
rect 299 3759 333 3775
rect 457 4751 491 4767
rect 457 3759 491 3775
rect 615 4751 649 4767
rect 615 3759 649 3775
rect 773 4751 807 4767
rect 773 3759 807 3775
rect 931 4751 965 4767
rect 931 3759 965 3775
rect 1089 4751 1123 4767
rect 1089 3759 1123 3775
rect 1247 4751 1281 4767
rect 1247 3759 1281 3775
rect 1405 4751 1439 4767
rect 1405 3759 1439 3775
rect 1563 4751 1597 4767
rect 1563 3759 1597 3775
rect -1551 3691 -1535 3725
rect -1467 3691 -1451 3725
rect -1393 3691 -1377 3725
rect -1309 3691 -1293 3725
rect -1235 3691 -1219 3725
rect -1151 3691 -1135 3725
rect -1077 3691 -1061 3725
rect -993 3691 -977 3725
rect -919 3691 -903 3725
rect -835 3691 -819 3725
rect -761 3691 -745 3725
rect -677 3691 -661 3725
rect -603 3691 -587 3725
rect -519 3691 -503 3725
rect -445 3691 -429 3725
rect -361 3691 -345 3725
rect -287 3691 -271 3725
rect -203 3691 -187 3725
rect -129 3691 -113 3725
rect -45 3691 -29 3725
rect 29 3691 45 3725
rect 113 3691 129 3725
rect 187 3691 203 3725
rect 271 3691 287 3725
rect 345 3691 361 3725
rect 429 3691 445 3725
rect 503 3691 519 3725
rect 587 3691 603 3725
rect 661 3691 677 3725
rect 745 3691 761 3725
rect 819 3691 835 3725
rect 903 3691 919 3725
rect 977 3691 993 3725
rect 1061 3691 1077 3725
rect 1135 3691 1151 3725
rect 1219 3691 1235 3725
rect 1293 3691 1309 3725
rect 1377 3691 1393 3725
rect 1451 3691 1467 3725
rect 1535 3691 1551 3725
rect -1551 3583 -1535 3617
rect -1467 3583 -1451 3617
rect -1393 3583 -1377 3617
rect -1309 3583 -1293 3617
rect -1235 3583 -1219 3617
rect -1151 3583 -1135 3617
rect -1077 3583 -1061 3617
rect -993 3583 -977 3617
rect -919 3583 -903 3617
rect -835 3583 -819 3617
rect -761 3583 -745 3617
rect -677 3583 -661 3617
rect -603 3583 -587 3617
rect -519 3583 -503 3617
rect -445 3583 -429 3617
rect -361 3583 -345 3617
rect -287 3583 -271 3617
rect -203 3583 -187 3617
rect -129 3583 -113 3617
rect -45 3583 -29 3617
rect 29 3583 45 3617
rect 113 3583 129 3617
rect 187 3583 203 3617
rect 271 3583 287 3617
rect 345 3583 361 3617
rect 429 3583 445 3617
rect 503 3583 519 3617
rect 587 3583 603 3617
rect 661 3583 677 3617
rect 745 3583 761 3617
rect 819 3583 835 3617
rect 903 3583 919 3617
rect 977 3583 993 3617
rect 1061 3583 1077 3617
rect 1135 3583 1151 3617
rect 1219 3583 1235 3617
rect 1293 3583 1309 3617
rect 1377 3583 1393 3617
rect 1451 3583 1467 3617
rect 1535 3583 1551 3617
rect -1597 3533 -1563 3549
rect -1597 2541 -1563 2557
rect -1439 3533 -1405 3549
rect -1439 2541 -1405 2557
rect -1281 3533 -1247 3549
rect -1281 2541 -1247 2557
rect -1123 3533 -1089 3549
rect -1123 2541 -1089 2557
rect -965 3533 -931 3549
rect -965 2541 -931 2557
rect -807 3533 -773 3549
rect -807 2541 -773 2557
rect -649 3533 -615 3549
rect -649 2541 -615 2557
rect -491 3533 -457 3549
rect -491 2541 -457 2557
rect -333 3533 -299 3549
rect -333 2541 -299 2557
rect -175 3533 -141 3549
rect -175 2541 -141 2557
rect -17 3533 17 3549
rect -17 2541 17 2557
rect 141 3533 175 3549
rect 141 2541 175 2557
rect 299 3533 333 3549
rect 299 2541 333 2557
rect 457 3533 491 3549
rect 457 2541 491 2557
rect 615 3533 649 3549
rect 615 2541 649 2557
rect 773 3533 807 3549
rect 773 2541 807 2557
rect 931 3533 965 3549
rect 931 2541 965 2557
rect 1089 3533 1123 3549
rect 1089 2541 1123 2557
rect 1247 3533 1281 3549
rect 1247 2541 1281 2557
rect 1405 3533 1439 3549
rect 1405 2541 1439 2557
rect 1563 3533 1597 3549
rect 1563 2541 1597 2557
rect -1551 2473 -1535 2507
rect -1467 2473 -1451 2507
rect -1393 2473 -1377 2507
rect -1309 2473 -1293 2507
rect -1235 2473 -1219 2507
rect -1151 2473 -1135 2507
rect -1077 2473 -1061 2507
rect -993 2473 -977 2507
rect -919 2473 -903 2507
rect -835 2473 -819 2507
rect -761 2473 -745 2507
rect -677 2473 -661 2507
rect -603 2473 -587 2507
rect -519 2473 -503 2507
rect -445 2473 -429 2507
rect -361 2473 -345 2507
rect -287 2473 -271 2507
rect -203 2473 -187 2507
rect -129 2473 -113 2507
rect -45 2473 -29 2507
rect 29 2473 45 2507
rect 113 2473 129 2507
rect 187 2473 203 2507
rect 271 2473 287 2507
rect 345 2473 361 2507
rect 429 2473 445 2507
rect 503 2473 519 2507
rect 587 2473 603 2507
rect 661 2473 677 2507
rect 745 2473 761 2507
rect 819 2473 835 2507
rect 903 2473 919 2507
rect 977 2473 993 2507
rect 1061 2473 1077 2507
rect 1135 2473 1151 2507
rect 1219 2473 1235 2507
rect 1293 2473 1309 2507
rect 1377 2473 1393 2507
rect 1451 2473 1467 2507
rect 1535 2473 1551 2507
rect -1551 2365 -1535 2399
rect -1467 2365 -1451 2399
rect -1393 2365 -1377 2399
rect -1309 2365 -1293 2399
rect -1235 2365 -1219 2399
rect -1151 2365 -1135 2399
rect -1077 2365 -1061 2399
rect -993 2365 -977 2399
rect -919 2365 -903 2399
rect -835 2365 -819 2399
rect -761 2365 -745 2399
rect -677 2365 -661 2399
rect -603 2365 -587 2399
rect -519 2365 -503 2399
rect -445 2365 -429 2399
rect -361 2365 -345 2399
rect -287 2365 -271 2399
rect -203 2365 -187 2399
rect -129 2365 -113 2399
rect -45 2365 -29 2399
rect 29 2365 45 2399
rect 113 2365 129 2399
rect 187 2365 203 2399
rect 271 2365 287 2399
rect 345 2365 361 2399
rect 429 2365 445 2399
rect 503 2365 519 2399
rect 587 2365 603 2399
rect 661 2365 677 2399
rect 745 2365 761 2399
rect 819 2365 835 2399
rect 903 2365 919 2399
rect 977 2365 993 2399
rect 1061 2365 1077 2399
rect 1135 2365 1151 2399
rect 1219 2365 1235 2399
rect 1293 2365 1309 2399
rect 1377 2365 1393 2399
rect 1451 2365 1467 2399
rect 1535 2365 1551 2399
rect -1597 2315 -1563 2331
rect -1597 1323 -1563 1339
rect -1439 2315 -1405 2331
rect -1439 1323 -1405 1339
rect -1281 2315 -1247 2331
rect -1281 1323 -1247 1339
rect -1123 2315 -1089 2331
rect -1123 1323 -1089 1339
rect -965 2315 -931 2331
rect -965 1323 -931 1339
rect -807 2315 -773 2331
rect -807 1323 -773 1339
rect -649 2315 -615 2331
rect -649 1323 -615 1339
rect -491 2315 -457 2331
rect -491 1323 -457 1339
rect -333 2315 -299 2331
rect -333 1323 -299 1339
rect -175 2315 -141 2331
rect -175 1323 -141 1339
rect -17 2315 17 2331
rect -17 1323 17 1339
rect 141 2315 175 2331
rect 141 1323 175 1339
rect 299 2315 333 2331
rect 299 1323 333 1339
rect 457 2315 491 2331
rect 457 1323 491 1339
rect 615 2315 649 2331
rect 615 1323 649 1339
rect 773 2315 807 2331
rect 773 1323 807 1339
rect 931 2315 965 2331
rect 931 1323 965 1339
rect 1089 2315 1123 2331
rect 1089 1323 1123 1339
rect 1247 2315 1281 2331
rect 1247 1323 1281 1339
rect 1405 2315 1439 2331
rect 1405 1323 1439 1339
rect 1563 2315 1597 2331
rect 1563 1323 1597 1339
rect -1551 1255 -1535 1289
rect -1467 1255 -1451 1289
rect -1393 1255 -1377 1289
rect -1309 1255 -1293 1289
rect -1235 1255 -1219 1289
rect -1151 1255 -1135 1289
rect -1077 1255 -1061 1289
rect -993 1255 -977 1289
rect -919 1255 -903 1289
rect -835 1255 -819 1289
rect -761 1255 -745 1289
rect -677 1255 -661 1289
rect -603 1255 -587 1289
rect -519 1255 -503 1289
rect -445 1255 -429 1289
rect -361 1255 -345 1289
rect -287 1255 -271 1289
rect -203 1255 -187 1289
rect -129 1255 -113 1289
rect -45 1255 -29 1289
rect 29 1255 45 1289
rect 113 1255 129 1289
rect 187 1255 203 1289
rect 271 1255 287 1289
rect 345 1255 361 1289
rect 429 1255 445 1289
rect 503 1255 519 1289
rect 587 1255 603 1289
rect 661 1255 677 1289
rect 745 1255 761 1289
rect 819 1255 835 1289
rect 903 1255 919 1289
rect 977 1255 993 1289
rect 1061 1255 1077 1289
rect 1135 1255 1151 1289
rect 1219 1255 1235 1289
rect 1293 1255 1309 1289
rect 1377 1255 1393 1289
rect 1451 1255 1467 1289
rect 1535 1255 1551 1289
rect -1551 1147 -1535 1181
rect -1467 1147 -1451 1181
rect -1393 1147 -1377 1181
rect -1309 1147 -1293 1181
rect -1235 1147 -1219 1181
rect -1151 1147 -1135 1181
rect -1077 1147 -1061 1181
rect -993 1147 -977 1181
rect -919 1147 -903 1181
rect -835 1147 -819 1181
rect -761 1147 -745 1181
rect -677 1147 -661 1181
rect -603 1147 -587 1181
rect -519 1147 -503 1181
rect -445 1147 -429 1181
rect -361 1147 -345 1181
rect -287 1147 -271 1181
rect -203 1147 -187 1181
rect -129 1147 -113 1181
rect -45 1147 -29 1181
rect 29 1147 45 1181
rect 113 1147 129 1181
rect 187 1147 203 1181
rect 271 1147 287 1181
rect 345 1147 361 1181
rect 429 1147 445 1181
rect 503 1147 519 1181
rect 587 1147 603 1181
rect 661 1147 677 1181
rect 745 1147 761 1181
rect 819 1147 835 1181
rect 903 1147 919 1181
rect 977 1147 993 1181
rect 1061 1147 1077 1181
rect 1135 1147 1151 1181
rect 1219 1147 1235 1181
rect 1293 1147 1309 1181
rect 1377 1147 1393 1181
rect 1451 1147 1467 1181
rect 1535 1147 1551 1181
rect -1597 1097 -1563 1113
rect -1597 105 -1563 121
rect -1439 1097 -1405 1113
rect -1439 105 -1405 121
rect -1281 1097 -1247 1113
rect -1281 105 -1247 121
rect -1123 1097 -1089 1113
rect -1123 105 -1089 121
rect -965 1097 -931 1113
rect -965 105 -931 121
rect -807 1097 -773 1113
rect -807 105 -773 121
rect -649 1097 -615 1113
rect -649 105 -615 121
rect -491 1097 -457 1113
rect -491 105 -457 121
rect -333 1097 -299 1113
rect -333 105 -299 121
rect -175 1097 -141 1113
rect -175 105 -141 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 141 1097 175 1113
rect 141 105 175 121
rect 299 1097 333 1113
rect 299 105 333 121
rect 457 1097 491 1113
rect 457 105 491 121
rect 615 1097 649 1113
rect 615 105 649 121
rect 773 1097 807 1113
rect 773 105 807 121
rect 931 1097 965 1113
rect 931 105 965 121
rect 1089 1097 1123 1113
rect 1089 105 1123 121
rect 1247 1097 1281 1113
rect 1247 105 1281 121
rect 1405 1097 1439 1113
rect 1405 105 1439 121
rect 1563 1097 1597 1113
rect 1563 105 1597 121
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect -1597 -121 -1563 -105
rect -1597 -1113 -1563 -1097
rect -1439 -121 -1405 -105
rect -1439 -1113 -1405 -1097
rect -1281 -121 -1247 -105
rect -1281 -1113 -1247 -1097
rect -1123 -121 -1089 -105
rect -1123 -1113 -1089 -1097
rect -965 -121 -931 -105
rect -965 -1113 -931 -1097
rect -807 -121 -773 -105
rect -807 -1113 -773 -1097
rect -649 -121 -615 -105
rect -649 -1113 -615 -1097
rect -491 -121 -457 -105
rect -491 -1113 -457 -1097
rect -333 -121 -299 -105
rect -333 -1113 -299 -1097
rect -175 -121 -141 -105
rect -175 -1113 -141 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 141 -121 175 -105
rect 141 -1113 175 -1097
rect 299 -121 333 -105
rect 299 -1113 333 -1097
rect 457 -121 491 -105
rect 457 -1113 491 -1097
rect 615 -121 649 -105
rect 615 -1113 649 -1097
rect 773 -121 807 -105
rect 773 -1113 807 -1097
rect 931 -121 965 -105
rect 931 -1113 965 -1097
rect 1089 -121 1123 -105
rect 1089 -1113 1123 -1097
rect 1247 -121 1281 -105
rect 1247 -1113 1281 -1097
rect 1405 -121 1439 -105
rect 1405 -1113 1439 -1097
rect 1563 -121 1597 -105
rect 1563 -1113 1597 -1097
rect -1551 -1181 -1535 -1147
rect -1467 -1181 -1451 -1147
rect -1393 -1181 -1377 -1147
rect -1309 -1181 -1293 -1147
rect -1235 -1181 -1219 -1147
rect -1151 -1181 -1135 -1147
rect -1077 -1181 -1061 -1147
rect -993 -1181 -977 -1147
rect -919 -1181 -903 -1147
rect -835 -1181 -819 -1147
rect -761 -1181 -745 -1147
rect -677 -1181 -661 -1147
rect -603 -1181 -587 -1147
rect -519 -1181 -503 -1147
rect -445 -1181 -429 -1147
rect -361 -1181 -345 -1147
rect -287 -1181 -271 -1147
rect -203 -1181 -187 -1147
rect -129 -1181 -113 -1147
rect -45 -1181 -29 -1147
rect 29 -1181 45 -1147
rect 113 -1181 129 -1147
rect 187 -1181 203 -1147
rect 271 -1181 287 -1147
rect 345 -1181 361 -1147
rect 429 -1181 445 -1147
rect 503 -1181 519 -1147
rect 587 -1181 603 -1147
rect 661 -1181 677 -1147
rect 745 -1181 761 -1147
rect 819 -1181 835 -1147
rect 903 -1181 919 -1147
rect 977 -1181 993 -1147
rect 1061 -1181 1077 -1147
rect 1135 -1181 1151 -1147
rect 1219 -1181 1235 -1147
rect 1293 -1181 1309 -1147
rect 1377 -1181 1393 -1147
rect 1451 -1181 1467 -1147
rect 1535 -1181 1551 -1147
rect -1551 -1289 -1535 -1255
rect -1467 -1289 -1451 -1255
rect -1393 -1289 -1377 -1255
rect -1309 -1289 -1293 -1255
rect -1235 -1289 -1219 -1255
rect -1151 -1289 -1135 -1255
rect -1077 -1289 -1061 -1255
rect -993 -1289 -977 -1255
rect -919 -1289 -903 -1255
rect -835 -1289 -819 -1255
rect -761 -1289 -745 -1255
rect -677 -1289 -661 -1255
rect -603 -1289 -587 -1255
rect -519 -1289 -503 -1255
rect -445 -1289 -429 -1255
rect -361 -1289 -345 -1255
rect -287 -1289 -271 -1255
rect -203 -1289 -187 -1255
rect -129 -1289 -113 -1255
rect -45 -1289 -29 -1255
rect 29 -1289 45 -1255
rect 113 -1289 129 -1255
rect 187 -1289 203 -1255
rect 271 -1289 287 -1255
rect 345 -1289 361 -1255
rect 429 -1289 445 -1255
rect 503 -1289 519 -1255
rect 587 -1289 603 -1255
rect 661 -1289 677 -1255
rect 745 -1289 761 -1255
rect 819 -1289 835 -1255
rect 903 -1289 919 -1255
rect 977 -1289 993 -1255
rect 1061 -1289 1077 -1255
rect 1135 -1289 1151 -1255
rect 1219 -1289 1235 -1255
rect 1293 -1289 1309 -1255
rect 1377 -1289 1393 -1255
rect 1451 -1289 1467 -1255
rect 1535 -1289 1551 -1255
rect -1597 -1339 -1563 -1323
rect -1597 -2331 -1563 -2315
rect -1439 -1339 -1405 -1323
rect -1439 -2331 -1405 -2315
rect -1281 -1339 -1247 -1323
rect -1281 -2331 -1247 -2315
rect -1123 -1339 -1089 -1323
rect -1123 -2331 -1089 -2315
rect -965 -1339 -931 -1323
rect -965 -2331 -931 -2315
rect -807 -1339 -773 -1323
rect -807 -2331 -773 -2315
rect -649 -1339 -615 -1323
rect -649 -2331 -615 -2315
rect -491 -1339 -457 -1323
rect -491 -2331 -457 -2315
rect -333 -1339 -299 -1323
rect -333 -2331 -299 -2315
rect -175 -1339 -141 -1323
rect -175 -2331 -141 -2315
rect -17 -1339 17 -1323
rect -17 -2331 17 -2315
rect 141 -1339 175 -1323
rect 141 -2331 175 -2315
rect 299 -1339 333 -1323
rect 299 -2331 333 -2315
rect 457 -1339 491 -1323
rect 457 -2331 491 -2315
rect 615 -1339 649 -1323
rect 615 -2331 649 -2315
rect 773 -1339 807 -1323
rect 773 -2331 807 -2315
rect 931 -1339 965 -1323
rect 931 -2331 965 -2315
rect 1089 -1339 1123 -1323
rect 1089 -2331 1123 -2315
rect 1247 -1339 1281 -1323
rect 1247 -2331 1281 -2315
rect 1405 -1339 1439 -1323
rect 1405 -2331 1439 -2315
rect 1563 -1339 1597 -1323
rect 1563 -2331 1597 -2315
rect -1551 -2399 -1535 -2365
rect -1467 -2399 -1451 -2365
rect -1393 -2399 -1377 -2365
rect -1309 -2399 -1293 -2365
rect -1235 -2399 -1219 -2365
rect -1151 -2399 -1135 -2365
rect -1077 -2399 -1061 -2365
rect -993 -2399 -977 -2365
rect -919 -2399 -903 -2365
rect -835 -2399 -819 -2365
rect -761 -2399 -745 -2365
rect -677 -2399 -661 -2365
rect -603 -2399 -587 -2365
rect -519 -2399 -503 -2365
rect -445 -2399 -429 -2365
rect -361 -2399 -345 -2365
rect -287 -2399 -271 -2365
rect -203 -2399 -187 -2365
rect -129 -2399 -113 -2365
rect -45 -2399 -29 -2365
rect 29 -2399 45 -2365
rect 113 -2399 129 -2365
rect 187 -2399 203 -2365
rect 271 -2399 287 -2365
rect 345 -2399 361 -2365
rect 429 -2399 445 -2365
rect 503 -2399 519 -2365
rect 587 -2399 603 -2365
rect 661 -2399 677 -2365
rect 745 -2399 761 -2365
rect 819 -2399 835 -2365
rect 903 -2399 919 -2365
rect 977 -2399 993 -2365
rect 1061 -2399 1077 -2365
rect 1135 -2399 1151 -2365
rect 1219 -2399 1235 -2365
rect 1293 -2399 1309 -2365
rect 1377 -2399 1393 -2365
rect 1451 -2399 1467 -2365
rect 1535 -2399 1551 -2365
rect -1551 -2507 -1535 -2473
rect -1467 -2507 -1451 -2473
rect -1393 -2507 -1377 -2473
rect -1309 -2507 -1293 -2473
rect -1235 -2507 -1219 -2473
rect -1151 -2507 -1135 -2473
rect -1077 -2507 -1061 -2473
rect -993 -2507 -977 -2473
rect -919 -2507 -903 -2473
rect -835 -2507 -819 -2473
rect -761 -2507 -745 -2473
rect -677 -2507 -661 -2473
rect -603 -2507 -587 -2473
rect -519 -2507 -503 -2473
rect -445 -2507 -429 -2473
rect -361 -2507 -345 -2473
rect -287 -2507 -271 -2473
rect -203 -2507 -187 -2473
rect -129 -2507 -113 -2473
rect -45 -2507 -29 -2473
rect 29 -2507 45 -2473
rect 113 -2507 129 -2473
rect 187 -2507 203 -2473
rect 271 -2507 287 -2473
rect 345 -2507 361 -2473
rect 429 -2507 445 -2473
rect 503 -2507 519 -2473
rect 587 -2507 603 -2473
rect 661 -2507 677 -2473
rect 745 -2507 761 -2473
rect 819 -2507 835 -2473
rect 903 -2507 919 -2473
rect 977 -2507 993 -2473
rect 1061 -2507 1077 -2473
rect 1135 -2507 1151 -2473
rect 1219 -2507 1235 -2473
rect 1293 -2507 1309 -2473
rect 1377 -2507 1393 -2473
rect 1451 -2507 1467 -2473
rect 1535 -2507 1551 -2473
rect -1597 -2557 -1563 -2541
rect -1597 -3549 -1563 -3533
rect -1439 -2557 -1405 -2541
rect -1439 -3549 -1405 -3533
rect -1281 -2557 -1247 -2541
rect -1281 -3549 -1247 -3533
rect -1123 -2557 -1089 -2541
rect -1123 -3549 -1089 -3533
rect -965 -2557 -931 -2541
rect -965 -3549 -931 -3533
rect -807 -2557 -773 -2541
rect -807 -3549 -773 -3533
rect -649 -2557 -615 -2541
rect -649 -3549 -615 -3533
rect -491 -2557 -457 -2541
rect -491 -3549 -457 -3533
rect -333 -2557 -299 -2541
rect -333 -3549 -299 -3533
rect -175 -2557 -141 -2541
rect -175 -3549 -141 -3533
rect -17 -2557 17 -2541
rect -17 -3549 17 -3533
rect 141 -2557 175 -2541
rect 141 -3549 175 -3533
rect 299 -2557 333 -2541
rect 299 -3549 333 -3533
rect 457 -2557 491 -2541
rect 457 -3549 491 -3533
rect 615 -2557 649 -2541
rect 615 -3549 649 -3533
rect 773 -2557 807 -2541
rect 773 -3549 807 -3533
rect 931 -2557 965 -2541
rect 931 -3549 965 -3533
rect 1089 -2557 1123 -2541
rect 1089 -3549 1123 -3533
rect 1247 -2557 1281 -2541
rect 1247 -3549 1281 -3533
rect 1405 -2557 1439 -2541
rect 1405 -3549 1439 -3533
rect 1563 -2557 1597 -2541
rect 1563 -3549 1597 -3533
rect -1551 -3617 -1535 -3583
rect -1467 -3617 -1451 -3583
rect -1393 -3617 -1377 -3583
rect -1309 -3617 -1293 -3583
rect -1235 -3617 -1219 -3583
rect -1151 -3617 -1135 -3583
rect -1077 -3617 -1061 -3583
rect -993 -3617 -977 -3583
rect -919 -3617 -903 -3583
rect -835 -3617 -819 -3583
rect -761 -3617 -745 -3583
rect -677 -3617 -661 -3583
rect -603 -3617 -587 -3583
rect -519 -3617 -503 -3583
rect -445 -3617 -429 -3583
rect -361 -3617 -345 -3583
rect -287 -3617 -271 -3583
rect -203 -3617 -187 -3583
rect -129 -3617 -113 -3583
rect -45 -3617 -29 -3583
rect 29 -3617 45 -3583
rect 113 -3617 129 -3583
rect 187 -3617 203 -3583
rect 271 -3617 287 -3583
rect 345 -3617 361 -3583
rect 429 -3617 445 -3583
rect 503 -3617 519 -3583
rect 587 -3617 603 -3583
rect 661 -3617 677 -3583
rect 745 -3617 761 -3583
rect 819 -3617 835 -3583
rect 903 -3617 919 -3583
rect 977 -3617 993 -3583
rect 1061 -3617 1077 -3583
rect 1135 -3617 1151 -3583
rect 1219 -3617 1235 -3583
rect 1293 -3617 1309 -3583
rect 1377 -3617 1393 -3583
rect 1451 -3617 1467 -3583
rect 1535 -3617 1551 -3583
rect -1551 -3725 -1535 -3691
rect -1467 -3725 -1451 -3691
rect -1393 -3725 -1377 -3691
rect -1309 -3725 -1293 -3691
rect -1235 -3725 -1219 -3691
rect -1151 -3725 -1135 -3691
rect -1077 -3725 -1061 -3691
rect -993 -3725 -977 -3691
rect -919 -3725 -903 -3691
rect -835 -3725 -819 -3691
rect -761 -3725 -745 -3691
rect -677 -3725 -661 -3691
rect -603 -3725 -587 -3691
rect -519 -3725 -503 -3691
rect -445 -3725 -429 -3691
rect -361 -3725 -345 -3691
rect -287 -3725 -271 -3691
rect -203 -3725 -187 -3691
rect -129 -3725 -113 -3691
rect -45 -3725 -29 -3691
rect 29 -3725 45 -3691
rect 113 -3725 129 -3691
rect 187 -3725 203 -3691
rect 271 -3725 287 -3691
rect 345 -3725 361 -3691
rect 429 -3725 445 -3691
rect 503 -3725 519 -3691
rect 587 -3725 603 -3691
rect 661 -3725 677 -3691
rect 745 -3725 761 -3691
rect 819 -3725 835 -3691
rect 903 -3725 919 -3691
rect 977 -3725 993 -3691
rect 1061 -3725 1077 -3691
rect 1135 -3725 1151 -3691
rect 1219 -3725 1235 -3691
rect 1293 -3725 1309 -3691
rect 1377 -3725 1393 -3691
rect 1451 -3725 1467 -3691
rect 1535 -3725 1551 -3691
rect -1597 -3775 -1563 -3759
rect -1597 -4767 -1563 -4751
rect -1439 -3775 -1405 -3759
rect -1439 -4767 -1405 -4751
rect -1281 -3775 -1247 -3759
rect -1281 -4767 -1247 -4751
rect -1123 -3775 -1089 -3759
rect -1123 -4767 -1089 -4751
rect -965 -3775 -931 -3759
rect -965 -4767 -931 -4751
rect -807 -3775 -773 -3759
rect -807 -4767 -773 -4751
rect -649 -3775 -615 -3759
rect -649 -4767 -615 -4751
rect -491 -3775 -457 -3759
rect -491 -4767 -457 -4751
rect -333 -3775 -299 -3759
rect -333 -4767 -299 -4751
rect -175 -3775 -141 -3759
rect -175 -4767 -141 -4751
rect -17 -3775 17 -3759
rect -17 -4767 17 -4751
rect 141 -3775 175 -3759
rect 141 -4767 175 -4751
rect 299 -3775 333 -3759
rect 299 -4767 333 -4751
rect 457 -3775 491 -3759
rect 457 -4767 491 -4751
rect 615 -3775 649 -3759
rect 615 -4767 649 -4751
rect 773 -3775 807 -3759
rect 773 -4767 807 -4751
rect 931 -3775 965 -3759
rect 931 -4767 965 -4751
rect 1089 -3775 1123 -3759
rect 1089 -4767 1123 -4751
rect 1247 -3775 1281 -3759
rect 1247 -4767 1281 -4751
rect 1405 -3775 1439 -3759
rect 1405 -4767 1439 -4751
rect 1563 -3775 1597 -3759
rect 1563 -4767 1597 -4751
rect -1551 -4835 -1535 -4801
rect -1467 -4835 -1451 -4801
rect -1393 -4835 -1377 -4801
rect -1309 -4835 -1293 -4801
rect -1235 -4835 -1219 -4801
rect -1151 -4835 -1135 -4801
rect -1077 -4835 -1061 -4801
rect -993 -4835 -977 -4801
rect -919 -4835 -903 -4801
rect -835 -4835 -819 -4801
rect -761 -4835 -745 -4801
rect -677 -4835 -661 -4801
rect -603 -4835 -587 -4801
rect -519 -4835 -503 -4801
rect -445 -4835 -429 -4801
rect -361 -4835 -345 -4801
rect -287 -4835 -271 -4801
rect -203 -4835 -187 -4801
rect -129 -4835 -113 -4801
rect -45 -4835 -29 -4801
rect 29 -4835 45 -4801
rect 113 -4835 129 -4801
rect 187 -4835 203 -4801
rect 271 -4835 287 -4801
rect 345 -4835 361 -4801
rect 429 -4835 445 -4801
rect 503 -4835 519 -4801
rect 587 -4835 603 -4801
rect 661 -4835 677 -4801
rect 745 -4835 761 -4801
rect 819 -4835 835 -4801
rect 903 -4835 919 -4801
rect 977 -4835 993 -4801
rect 1061 -4835 1077 -4801
rect 1135 -4835 1151 -4801
rect 1219 -4835 1235 -4801
rect 1293 -4835 1309 -4801
rect 1377 -4835 1393 -4801
rect 1451 -4835 1467 -4801
rect 1535 -4835 1551 -4801
rect -1551 -4943 -1535 -4909
rect -1467 -4943 -1451 -4909
rect -1393 -4943 -1377 -4909
rect -1309 -4943 -1293 -4909
rect -1235 -4943 -1219 -4909
rect -1151 -4943 -1135 -4909
rect -1077 -4943 -1061 -4909
rect -993 -4943 -977 -4909
rect -919 -4943 -903 -4909
rect -835 -4943 -819 -4909
rect -761 -4943 -745 -4909
rect -677 -4943 -661 -4909
rect -603 -4943 -587 -4909
rect -519 -4943 -503 -4909
rect -445 -4943 -429 -4909
rect -361 -4943 -345 -4909
rect -287 -4943 -271 -4909
rect -203 -4943 -187 -4909
rect -129 -4943 -113 -4909
rect -45 -4943 -29 -4909
rect 29 -4943 45 -4909
rect 113 -4943 129 -4909
rect 187 -4943 203 -4909
rect 271 -4943 287 -4909
rect 345 -4943 361 -4909
rect 429 -4943 445 -4909
rect 503 -4943 519 -4909
rect 587 -4943 603 -4909
rect 661 -4943 677 -4909
rect 745 -4943 761 -4909
rect 819 -4943 835 -4909
rect 903 -4943 919 -4909
rect 977 -4943 993 -4909
rect 1061 -4943 1077 -4909
rect 1135 -4943 1151 -4909
rect 1219 -4943 1235 -4909
rect 1293 -4943 1309 -4909
rect 1377 -4943 1393 -4909
rect 1451 -4943 1467 -4909
rect 1535 -4943 1551 -4909
rect -1597 -4993 -1563 -4977
rect -1597 -5985 -1563 -5969
rect -1439 -4993 -1405 -4977
rect -1439 -5985 -1405 -5969
rect -1281 -4993 -1247 -4977
rect -1281 -5985 -1247 -5969
rect -1123 -4993 -1089 -4977
rect -1123 -5985 -1089 -5969
rect -965 -4993 -931 -4977
rect -965 -5985 -931 -5969
rect -807 -4993 -773 -4977
rect -807 -5985 -773 -5969
rect -649 -4993 -615 -4977
rect -649 -5985 -615 -5969
rect -491 -4993 -457 -4977
rect -491 -5985 -457 -5969
rect -333 -4993 -299 -4977
rect -333 -5985 -299 -5969
rect -175 -4993 -141 -4977
rect -175 -5985 -141 -5969
rect -17 -4993 17 -4977
rect -17 -5985 17 -5969
rect 141 -4993 175 -4977
rect 141 -5985 175 -5969
rect 299 -4993 333 -4977
rect 299 -5985 333 -5969
rect 457 -4993 491 -4977
rect 457 -5985 491 -5969
rect 615 -4993 649 -4977
rect 615 -5985 649 -5969
rect 773 -4993 807 -4977
rect 773 -5985 807 -5969
rect 931 -4993 965 -4977
rect 931 -5985 965 -5969
rect 1089 -4993 1123 -4977
rect 1089 -5985 1123 -5969
rect 1247 -4993 1281 -4977
rect 1247 -5985 1281 -5969
rect 1405 -4993 1439 -4977
rect 1405 -5985 1439 -5969
rect 1563 -4993 1597 -4977
rect 1563 -5985 1597 -5969
rect -1551 -6053 -1535 -6019
rect -1467 -6053 -1451 -6019
rect -1393 -6053 -1377 -6019
rect -1309 -6053 -1293 -6019
rect -1235 -6053 -1219 -6019
rect -1151 -6053 -1135 -6019
rect -1077 -6053 -1061 -6019
rect -993 -6053 -977 -6019
rect -919 -6053 -903 -6019
rect -835 -6053 -819 -6019
rect -761 -6053 -745 -6019
rect -677 -6053 -661 -6019
rect -603 -6053 -587 -6019
rect -519 -6053 -503 -6019
rect -445 -6053 -429 -6019
rect -361 -6053 -345 -6019
rect -287 -6053 -271 -6019
rect -203 -6053 -187 -6019
rect -129 -6053 -113 -6019
rect -45 -6053 -29 -6019
rect 29 -6053 45 -6019
rect 113 -6053 129 -6019
rect 187 -6053 203 -6019
rect 271 -6053 287 -6019
rect 345 -6053 361 -6019
rect 429 -6053 445 -6019
rect 503 -6053 519 -6019
rect 587 -6053 603 -6019
rect 661 -6053 677 -6019
rect 745 -6053 761 -6019
rect 819 -6053 835 -6019
rect 903 -6053 919 -6019
rect 977 -6053 993 -6019
rect 1061 -6053 1077 -6019
rect 1135 -6053 1151 -6019
rect 1219 -6053 1235 -6019
rect 1293 -6053 1309 -6019
rect 1377 -6053 1393 -6019
rect 1451 -6053 1467 -6019
rect 1535 -6053 1551 -6019
rect -1741 -6157 -1707 -6095
rect 1707 -6157 1741 -6095
rect -1741 -6191 -1645 -6157
rect 1645 -6191 1741 -6157
<< viali >>
rect -1535 6019 -1467 6053
rect -1377 6019 -1309 6053
rect -1219 6019 -1151 6053
rect -1061 6019 -993 6053
rect -903 6019 -835 6053
rect -745 6019 -677 6053
rect -587 6019 -519 6053
rect -429 6019 -361 6053
rect -271 6019 -203 6053
rect -113 6019 -45 6053
rect 45 6019 113 6053
rect 203 6019 271 6053
rect 361 6019 429 6053
rect 519 6019 587 6053
rect 677 6019 745 6053
rect 835 6019 903 6053
rect 993 6019 1061 6053
rect 1151 6019 1219 6053
rect 1309 6019 1377 6053
rect 1467 6019 1535 6053
rect -1597 4993 -1563 5969
rect -1439 4993 -1405 5969
rect -1281 4993 -1247 5969
rect -1123 4993 -1089 5969
rect -965 4993 -931 5969
rect -807 4993 -773 5969
rect -649 4993 -615 5969
rect -491 4993 -457 5969
rect -333 4993 -299 5969
rect -175 4993 -141 5969
rect -17 4993 17 5969
rect 141 4993 175 5969
rect 299 4993 333 5969
rect 457 4993 491 5969
rect 615 4993 649 5969
rect 773 4993 807 5969
rect 931 4993 965 5969
rect 1089 4993 1123 5969
rect 1247 4993 1281 5969
rect 1405 4993 1439 5969
rect 1563 4993 1597 5969
rect -1535 4909 -1467 4943
rect -1377 4909 -1309 4943
rect -1219 4909 -1151 4943
rect -1061 4909 -993 4943
rect -903 4909 -835 4943
rect -745 4909 -677 4943
rect -587 4909 -519 4943
rect -429 4909 -361 4943
rect -271 4909 -203 4943
rect -113 4909 -45 4943
rect 45 4909 113 4943
rect 203 4909 271 4943
rect 361 4909 429 4943
rect 519 4909 587 4943
rect 677 4909 745 4943
rect 835 4909 903 4943
rect 993 4909 1061 4943
rect 1151 4909 1219 4943
rect 1309 4909 1377 4943
rect 1467 4909 1535 4943
rect -1535 4801 -1467 4835
rect -1377 4801 -1309 4835
rect -1219 4801 -1151 4835
rect -1061 4801 -993 4835
rect -903 4801 -835 4835
rect -745 4801 -677 4835
rect -587 4801 -519 4835
rect -429 4801 -361 4835
rect -271 4801 -203 4835
rect -113 4801 -45 4835
rect 45 4801 113 4835
rect 203 4801 271 4835
rect 361 4801 429 4835
rect 519 4801 587 4835
rect 677 4801 745 4835
rect 835 4801 903 4835
rect 993 4801 1061 4835
rect 1151 4801 1219 4835
rect 1309 4801 1377 4835
rect 1467 4801 1535 4835
rect -1597 3775 -1563 4751
rect -1439 3775 -1405 4751
rect -1281 3775 -1247 4751
rect -1123 3775 -1089 4751
rect -965 3775 -931 4751
rect -807 3775 -773 4751
rect -649 3775 -615 4751
rect -491 3775 -457 4751
rect -333 3775 -299 4751
rect -175 3775 -141 4751
rect -17 3775 17 4751
rect 141 3775 175 4751
rect 299 3775 333 4751
rect 457 3775 491 4751
rect 615 3775 649 4751
rect 773 3775 807 4751
rect 931 3775 965 4751
rect 1089 3775 1123 4751
rect 1247 3775 1281 4751
rect 1405 3775 1439 4751
rect 1563 3775 1597 4751
rect -1535 3691 -1467 3725
rect -1377 3691 -1309 3725
rect -1219 3691 -1151 3725
rect -1061 3691 -993 3725
rect -903 3691 -835 3725
rect -745 3691 -677 3725
rect -587 3691 -519 3725
rect -429 3691 -361 3725
rect -271 3691 -203 3725
rect -113 3691 -45 3725
rect 45 3691 113 3725
rect 203 3691 271 3725
rect 361 3691 429 3725
rect 519 3691 587 3725
rect 677 3691 745 3725
rect 835 3691 903 3725
rect 993 3691 1061 3725
rect 1151 3691 1219 3725
rect 1309 3691 1377 3725
rect 1467 3691 1535 3725
rect -1535 3583 -1467 3617
rect -1377 3583 -1309 3617
rect -1219 3583 -1151 3617
rect -1061 3583 -993 3617
rect -903 3583 -835 3617
rect -745 3583 -677 3617
rect -587 3583 -519 3617
rect -429 3583 -361 3617
rect -271 3583 -203 3617
rect -113 3583 -45 3617
rect 45 3583 113 3617
rect 203 3583 271 3617
rect 361 3583 429 3617
rect 519 3583 587 3617
rect 677 3583 745 3617
rect 835 3583 903 3617
rect 993 3583 1061 3617
rect 1151 3583 1219 3617
rect 1309 3583 1377 3617
rect 1467 3583 1535 3617
rect -1597 2557 -1563 3533
rect -1439 2557 -1405 3533
rect -1281 2557 -1247 3533
rect -1123 2557 -1089 3533
rect -965 2557 -931 3533
rect -807 2557 -773 3533
rect -649 2557 -615 3533
rect -491 2557 -457 3533
rect -333 2557 -299 3533
rect -175 2557 -141 3533
rect -17 2557 17 3533
rect 141 2557 175 3533
rect 299 2557 333 3533
rect 457 2557 491 3533
rect 615 2557 649 3533
rect 773 2557 807 3533
rect 931 2557 965 3533
rect 1089 2557 1123 3533
rect 1247 2557 1281 3533
rect 1405 2557 1439 3533
rect 1563 2557 1597 3533
rect -1535 2473 -1467 2507
rect -1377 2473 -1309 2507
rect -1219 2473 -1151 2507
rect -1061 2473 -993 2507
rect -903 2473 -835 2507
rect -745 2473 -677 2507
rect -587 2473 -519 2507
rect -429 2473 -361 2507
rect -271 2473 -203 2507
rect -113 2473 -45 2507
rect 45 2473 113 2507
rect 203 2473 271 2507
rect 361 2473 429 2507
rect 519 2473 587 2507
rect 677 2473 745 2507
rect 835 2473 903 2507
rect 993 2473 1061 2507
rect 1151 2473 1219 2507
rect 1309 2473 1377 2507
rect 1467 2473 1535 2507
rect -1535 2365 -1467 2399
rect -1377 2365 -1309 2399
rect -1219 2365 -1151 2399
rect -1061 2365 -993 2399
rect -903 2365 -835 2399
rect -745 2365 -677 2399
rect -587 2365 -519 2399
rect -429 2365 -361 2399
rect -271 2365 -203 2399
rect -113 2365 -45 2399
rect 45 2365 113 2399
rect 203 2365 271 2399
rect 361 2365 429 2399
rect 519 2365 587 2399
rect 677 2365 745 2399
rect 835 2365 903 2399
rect 993 2365 1061 2399
rect 1151 2365 1219 2399
rect 1309 2365 1377 2399
rect 1467 2365 1535 2399
rect -1597 1339 -1563 2315
rect -1439 1339 -1405 2315
rect -1281 1339 -1247 2315
rect -1123 1339 -1089 2315
rect -965 1339 -931 2315
rect -807 1339 -773 2315
rect -649 1339 -615 2315
rect -491 1339 -457 2315
rect -333 1339 -299 2315
rect -175 1339 -141 2315
rect -17 1339 17 2315
rect 141 1339 175 2315
rect 299 1339 333 2315
rect 457 1339 491 2315
rect 615 1339 649 2315
rect 773 1339 807 2315
rect 931 1339 965 2315
rect 1089 1339 1123 2315
rect 1247 1339 1281 2315
rect 1405 1339 1439 2315
rect 1563 1339 1597 2315
rect -1535 1255 -1467 1289
rect -1377 1255 -1309 1289
rect -1219 1255 -1151 1289
rect -1061 1255 -993 1289
rect -903 1255 -835 1289
rect -745 1255 -677 1289
rect -587 1255 -519 1289
rect -429 1255 -361 1289
rect -271 1255 -203 1289
rect -113 1255 -45 1289
rect 45 1255 113 1289
rect 203 1255 271 1289
rect 361 1255 429 1289
rect 519 1255 587 1289
rect 677 1255 745 1289
rect 835 1255 903 1289
rect 993 1255 1061 1289
rect 1151 1255 1219 1289
rect 1309 1255 1377 1289
rect 1467 1255 1535 1289
rect -1535 1147 -1467 1181
rect -1377 1147 -1309 1181
rect -1219 1147 -1151 1181
rect -1061 1147 -993 1181
rect -903 1147 -835 1181
rect -745 1147 -677 1181
rect -587 1147 -519 1181
rect -429 1147 -361 1181
rect -271 1147 -203 1181
rect -113 1147 -45 1181
rect 45 1147 113 1181
rect 203 1147 271 1181
rect 361 1147 429 1181
rect 519 1147 587 1181
rect 677 1147 745 1181
rect 835 1147 903 1181
rect 993 1147 1061 1181
rect 1151 1147 1219 1181
rect 1309 1147 1377 1181
rect 1467 1147 1535 1181
rect -1597 121 -1563 1097
rect -1439 121 -1405 1097
rect -1281 121 -1247 1097
rect -1123 121 -1089 1097
rect -965 121 -931 1097
rect -807 121 -773 1097
rect -649 121 -615 1097
rect -491 121 -457 1097
rect -333 121 -299 1097
rect -175 121 -141 1097
rect -17 121 17 1097
rect 141 121 175 1097
rect 299 121 333 1097
rect 457 121 491 1097
rect 615 121 649 1097
rect 773 121 807 1097
rect 931 121 965 1097
rect 1089 121 1123 1097
rect 1247 121 1281 1097
rect 1405 121 1439 1097
rect 1563 121 1597 1097
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect -1597 -1097 -1563 -121
rect -1439 -1097 -1405 -121
rect -1281 -1097 -1247 -121
rect -1123 -1097 -1089 -121
rect -965 -1097 -931 -121
rect -807 -1097 -773 -121
rect -649 -1097 -615 -121
rect -491 -1097 -457 -121
rect -333 -1097 -299 -121
rect -175 -1097 -141 -121
rect -17 -1097 17 -121
rect 141 -1097 175 -121
rect 299 -1097 333 -121
rect 457 -1097 491 -121
rect 615 -1097 649 -121
rect 773 -1097 807 -121
rect 931 -1097 965 -121
rect 1089 -1097 1123 -121
rect 1247 -1097 1281 -121
rect 1405 -1097 1439 -121
rect 1563 -1097 1597 -121
rect -1535 -1181 -1467 -1147
rect -1377 -1181 -1309 -1147
rect -1219 -1181 -1151 -1147
rect -1061 -1181 -993 -1147
rect -903 -1181 -835 -1147
rect -745 -1181 -677 -1147
rect -587 -1181 -519 -1147
rect -429 -1181 -361 -1147
rect -271 -1181 -203 -1147
rect -113 -1181 -45 -1147
rect 45 -1181 113 -1147
rect 203 -1181 271 -1147
rect 361 -1181 429 -1147
rect 519 -1181 587 -1147
rect 677 -1181 745 -1147
rect 835 -1181 903 -1147
rect 993 -1181 1061 -1147
rect 1151 -1181 1219 -1147
rect 1309 -1181 1377 -1147
rect 1467 -1181 1535 -1147
rect -1535 -1289 -1467 -1255
rect -1377 -1289 -1309 -1255
rect -1219 -1289 -1151 -1255
rect -1061 -1289 -993 -1255
rect -903 -1289 -835 -1255
rect -745 -1289 -677 -1255
rect -587 -1289 -519 -1255
rect -429 -1289 -361 -1255
rect -271 -1289 -203 -1255
rect -113 -1289 -45 -1255
rect 45 -1289 113 -1255
rect 203 -1289 271 -1255
rect 361 -1289 429 -1255
rect 519 -1289 587 -1255
rect 677 -1289 745 -1255
rect 835 -1289 903 -1255
rect 993 -1289 1061 -1255
rect 1151 -1289 1219 -1255
rect 1309 -1289 1377 -1255
rect 1467 -1289 1535 -1255
rect -1597 -2315 -1563 -1339
rect -1439 -2315 -1405 -1339
rect -1281 -2315 -1247 -1339
rect -1123 -2315 -1089 -1339
rect -965 -2315 -931 -1339
rect -807 -2315 -773 -1339
rect -649 -2315 -615 -1339
rect -491 -2315 -457 -1339
rect -333 -2315 -299 -1339
rect -175 -2315 -141 -1339
rect -17 -2315 17 -1339
rect 141 -2315 175 -1339
rect 299 -2315 333 -1339
rect 457 -2315 491 -1339
rect 615 -2315 649 -1339
rect 773 -2315 807 -1339
rect 931 -2315 965 -1339
rect 1089 -2315 1123 -1339
rect 1247 -2315 1281 -1339
rect 1405 -2315 1439 -1339
rect 1563 -2315 1597 -1339
rect -1535 -2399 -1467 -2365
rect -1377 -2399 -1309 -2365
rect -1219 -2399 -1151 -2365
rect -1061 -2399 -993 -2365
rect -903 -2399 -835 -2365
rect -745 -2399 -677 -2365
rect -587 -2399 -519 -2365
rect -429 -2399 -361 -2365
rect -271 -2399 -203 -2365
rect -113 -2399 -45 -2365
rect 45 -2399 113 -2365
rect 203 -2399 271 -2365
rect 361 -2399 429 -2365
rect 519 -2399 587 -2365
rect 677 -2399 745 -2365
rect 835 -2399 903 -2365
rect 993 -2399 1061 -2365
rect 1151 -2399 1219 -2365
rect 1309 -2399 1377 -2365
rect 1467 -2399 1535 -2365
rect -1535 -2507 -1467 -2473
rect -1377 -2507 -1309 -2473
rect -1219 -2507 -1151 -2473
rect -1061 -2507 -993 -2473
rect -903 -2507 -835 -2473
rect -745 -2507 -677 -2473
rect -587 -2507 -519 -2473
rect -429 -2507 -361 -2473
rect -271 -2507 -203 -2473
rect -113 -2507 -45 -2473
rect 45 -2507 113 -2473
rect 203 -2507 271 -2473
rect 361 -2507 429 -2473
rect 519 -2507 587 -2473
rect 677 -2507 745 -2473
rect 835 -2507 903 -2473
rect 993 -2507 1061 -2473
rect 1151 -2507 1219 -2473
rect 1309 -2507 1377 -2473
rect 1467 -2507 1535 -2473
rect -1597 -3533 -1563 -2557
rect -1439 -3533 -1405 -2557
rect -1281 -3533 -1247 -2557
rect -1123 -3533 -1089 -2557
rect -965 -3533 -931 -2557
rect -807 -3533 -773 -2557
rect -649 -3533 -615 -2557
rect -491 -3533 -457 -2557
rect -333 -3533 -299 -2557
rect -175 -3533 -141 -2557
rect -17 -3533 17 -2557
rect 141 -3533 175 -2557
rect 299 -3533 333 -2557
rect 457 -3533 491 -2557
rect 615 -3533 649 -2557
rect 773 -3533 807 -2557
rect 931 -3533 965 -2557
rect 1089 -3533 1123 -2557
rect 1247 -3533 1281 -2557
rect 1405 -3533 1439 -2557
rect 1563 -3533 1597 -2557
rect -1535 -3617 -1467 -3583
rect -1377 -3617 -1309 -3583
rect -1219 -3617 -1151 -3583
rect -1061 -3617 -993 -3583
rect -903 -3617 -835 -3583
rect -745 -3617 -677 -3583
rect -587 -3617 -519 -3583
rect -429 -3617 -361 -3583
rect -271 -3617 -203 -3583
rect -113 -3617 -45 -3583
rect 45 -3617 113 -3583
rect 203 -3617 271 -3583
rect 361 -3617 429 -3583
rect 519 -3617 587 -3583
rect 677 -3617 745 -3583
rect 835 -3617 903 -3583
rect 993 -3617 1061 -3583
rect 1151 -3617 1219 -3583
rect 1309 -3617 1377 -3583
rect 1467 -3617 1535 -3583
rect -1535 -3725 -1467 -3691
rect -1377 -3725 -1309 -3691
rect -1219 -3725 -1151 -3691
rect -1061 -3725 -993 -3691
rect -903 -3725 -835 -3691
rect -745 -3725 -677 -3691
rect -587 -3725 -519 -3691
rect -429 -3725 -361 -3691
rect -271 -3725 -203 -3691
rect -113 -3725 -45 -3691
rect 45 -3725 113 -3691
rect 203 -3725 271 -3691
rect 361 -3725 429 -3691
rect 519 -3725 587 -3691
rect 677 -3725 745 -3691
rect 835 -3725 903 -3691
rect 993 -3725 1061 -3691
rect 1151 -3725 1219 -3691
rect 1309 -3725 1377 -3691
rect 1467 -3725 1535 -3691
rect -1597 -4751 -1563 -3775
rect -1439 -4751 -1405 -3775
rect -1281 -4751 -1247 -3775
rect -1123 -4751 -1089 -3775
rect -965 -4751 -931 -3775
rect -807 -4751 -773 -3775
rect -649 -4751 -615 -3775
rect -491 -4751 -457 -3775
rect -333 -4751 -299 -3775
rect -175 -4751 -141 -3775
rect -17 -4751 17 -3775
rect 141 -4751 175 -3775
rect 299 -4751 333 -3775
rect 457 -4751 491 -3775
rect 615 -4751 649 -3775
rect 773 -4751 807 -3775
rect 931 -4751 965 -3775
rect 1089 -4751 1123 -3775
rect 1247 -4751 1281 -3775
rect 1405 -4751 1439 -3775
rect 1563 -4751 1597 -3775
rect -1535 -4835 -1467 -4801
rect -1377 -4835 -1309 -4801
rect -1219 -4835 -1151 -4801
rect -1061 -4835 -993 -4801
rect -903 -4835 -835 -4801
rect -745 -4835 -677 -4801
rect -587 -4835 -519 -4801
rect -429 -4835 -361 -4801
rect -271 -4835 -203 -4801
rect -113 -4835 -45 -4801
rect 45 -4835 113 -4801
rect 203 -4835 271 -4801
rect 361 -4835 429 -4801
rect 519 -4835 587 -4801
rect 677 -4835 745 -4801
rect 835 -4835 903 -4801
rect 993 -4835 1061 -4801
rect 1151 -4835 1219 -4801
rect 1309 -4835 1377 -4801
rect 1467 -4835 1535 -4801
rect -1535 -4943 -1467 -4909
rect -1377 -4943 -1309 -4909
rect -1219 -4943 -1151 -4909
rect -1061 -4943 -993 -4909
rect -903 -4943 -835 -4909
rect -745 -4943 -677 -4909
rect -587 -4943 -519 -4909
rect -429 -4943 -361 -4909
rect -271 -4943 -203 -4909
rect -113 -4943 -45 -4909
rect 45 -4943 113 -4909
rect 203 -4943 271 -4909
rect 361 -4943 429 -4909
rect 519 -4943 587 -4909
rect 677 -4943 745 -4909
rect 835 -4943 903 -4909
rect 993 -4943 1061 -4909
rect 1151 -4943 1219 -4909
rect 1309 -4943 1377 -4909
rect 1467 -4943 1535 -4909
rect -1597 -5969 -1563 -4993
rect -1439 -5969 -1405 -4993
rect -1281 -5969 -1247 -4993
rect -1123 -5969 -1089 -4993
rect -965 -5969 -931 -4993
rect -807 -5969 -773 -4993
rect -649 -5969 -615 -4993
rect -491 -5969 -457 -4993
rect -333 -5969 -299 -4993
rect -175 -5969 -141 -4993
rect -17 -5969 17 -4993
rect 141 -5969 175 -4993
rect 299 -5969 333 -4993
rect 457 -5969 491 -4993
rect 615 -5969 649 -4993
rect 773 -5969 807 -4993
rect 931 -5969 965 -4993
rect 1089 -5969 1123 -4993
rect 1247 -5969 1281 -4993
rect 1405 -5969 1439 -4993
rect 1563 -5969 1597 -4993
rect -1535 -6053 -1467 -6019
rect -1377 -6053 -1309 -6019
rect -1219 -6053 -1151 -6019
rect -1061 -6053 -993 -6019
rect -903 -6053 -835 -6019
rect -745 -6053 -677 -6019
rect -587 -6053 -519 -6019
rect -429 -6053 -361 -6019
rect -271 -6053 -203 -6019
rect -113 -6053 -45 -6019
rect 45 -6053 113 -6019
rect 203 -6053 271 -6019
rect 361 -6053 429 -6019
rect 519 -6053 587 -6019
rect 677 -6053 745 -6019
rect 835 -6053 903 -6019
rect 993 -6053 1061 -6019
rect 1151 -6053 1219 -6019
rect 1309 -6053 1377 -6019
rect 1467 -6053 1535 -6019
<< metal1 >>
rect -1547 6053 -1455 6059
rect -1547 6019 -1535 6053
rect -1467 6019 -1455 6053
rect -1547 6013 -1455 6019
rect -1389 6053 -1297 6059
rect -1389 6019 -1377 6053
rect -1309 6019 -1297 6053
rect -1389 6013 -1297 6019
rect -1231 6053 -1139 6059
rect -1231 6019 -1219 6053
rect -1151 6019 -1139 6053
rect -1231 6013 -1139 6019
rect -1073 6053 -981 6059
rect -1073 6019 -1061 6053
rect -993 6019 -981 6053
rect -1073 6013 -981 6019
rect -915 6053 -823 6059
rect -915 6019 -903 6053
rect -835 6019 -823 6053
rect -915 6013 -823 6019
rect -757 6053 -665 6059
rect -757 6019 -745 6053
rect -677 6019 -665 6053
rect -757 6013 -665 6019
rect -599 6053 -507 6059
rect -599 6019 -587 6053
rect -519 6019 -507 6053
rect -599 6013 -507 6019
rect -441 6053 -349 6059
rect -441 6019 -429 6053
rect -361 6019 -349 6053
rect -441 6013 -349 6019
rect -283 6053 -191 6059
rect -283 6019 -271 6053
rect -203 6019 -191 6053
rect -283 6013 -191 6019
rect -125 6053 -33 6059
rect -125 6019 -113 6053
rect -45 6019 -33 6053
rect -125 6013 -33 6019
rect 33 6053 125 6059
rect 33 6019 45 6053
rect 113 6019 125 6053
rect 33 6013 125 6019
rect 191 6053 283 6059
rect 191 6019 203 6053
rect 271 6019 283 6053
rect 191 6013 283 6019
rect 349 6053 441 6059
rect 349 6019 361 6053
rect 429 6019 441 6053
rect 349 6013 441 6019
rect 507 6053 599 6059
rect 507 6019 519 6053
rect 587 6019 599 6053
rect 507 6013 599 6019
rect 665 6053 757 6059
rect 665 6019 677 6053
rect 745 6019 757 6053
rect 665 6013 757 6019
rect 823 6053 915 6059
rect 823 6019 835 6053
rect 903 6019 915 6053
rect 823 6013 915 6019
rect 981 6053 1073 6059
rect 981 6019 993 6053
rect 1061 6019 1073 6053
rect 981 6013 1073 6019
rect 1139 6053 1231 6059
rect 1139 6019 1151 6053
rect 1219 6019 1231 6053
rect 1139 6013 1231 6019
rect 1297 6053 1389 6059
rect 1297 6019 1309 6053
rect 1377 6019 1389 6053
rect 1297 6013 1389 6019
rect 1455 6053 1547 6059
rect 1455 6019 1467 6053
rect 1535 6019 1547 6053
rect 1455 6013 1547 6019
rect -1603 5969 -1557 5981
rect -1603 4993 -1597 5969
rect -1563 4993 -1557 5969
rect -1603 4981 -1557 4993
rect -1445 5969 -1399 5981
rect -1445 4993 -1439 5969
rect -1405 4993 -1399 5969
rect -1445 4981 -1399 4993
rect -1287 5969 -1241 5981
rect -1287 4993 -1281 5969
rect -1247 4993 -1241 5969
rect -1287 4981 -1241 4993
rect -1129 5969 -1083 5981
rect -1129 4993 -1123 5969
rect -1089 4993 -1083 5969
rect -1129 4981 -1083 4993
rect -971 5969 -925 5981
rect -971 4993 -965 5969
rect -931 4993 -925 5969
rect -971 4981 -925 4993
rect -813 5969 -767 5981
rect -813 4993 -807 5969
rect -773 4993 -767 5969
rect -813 4981 -767 4993
rect -655 5969 -609 5981
rect -655 4993 -649 5969
rect -615 4993 -609 5969
rect -655 4981 -609 4993
rect -497 5969 -451 5981
rect -497 4993 -491 5969
rect -457 4993 -451 5969
rect -497 4981 -451 4993
rect -339 5969 -293 5981
rect -339 4993 -333 5969
rect -299 4993 -293 5969
rect -339 4981 -293 4993
rect -181 5969 -135 5981
rect -181 4993 -175 5969
rect -141 4993 -135 5969
rect -181 4981 -135 4993
rect -23 5969 23 5981
rect -23 4993 -17 5969
rect 17 4993 23 5969
rect -23 4981 23 4993
rect 135 5969 181 5981
rect 135 4993 141 5969
rect 175 4993 181 5969
rect 135 4981 181 4993
rect 293 5969 339 5981
rect 293 4993 299 5969
rect 333 4993 339 5969
rect 293 4981 339 4993
rect 451 5969 497 5981
rect 451 4993 457 5969
rect 491 4993 497 5969
rect 451 4981 497 4993
rect 609 5969 655 5981
rect 609 4993 615 5969
rect 649 4993 655 5969
rect 609 4981 655 4993
rect 767 5969 813 5981
rect 767 4993 773 5969
rect 807 4993 813 5969
rect 767 4981 813 4993
rect 925 5969 971 5981
rect 925 4993 931 5969
rect 965 4993 971 5969
rect 925 4981 971 4993
rect 1083 5969 1129 5981
rect 1083 4993 1089 5969
rect 1123 4993 1129 5969
rect 1083 4981 1129 4993
rect 1241 5969 1287 5981
rect 1241 4993 1247 5969
rect 1281 4993 1287 5969
rect 1241 4981 1287 4993
rect 1399 5969 1445 5981
rect 1399 4993 1405 5969
rect 1439 4993 1445 5969
rect 1399 4981 1445 4993
rect 1557 5969 1603 5981
rect 1557 4993 1563 5969
rect 1597 4993 1603 5969
rect 1557 4981 1603 4993
rect -1547 4943 -1455 4949
rect -1547 4909 -1535 4943
rect -1467 4909 -1455 4943
rect -1547 4903 -1455 4909
rect -1389 4943 -1297 4949
rect -1389 4909 -1377 4943
rect -1309 4909 -1297 4943
rect -1389 4903 -1297 4909
rect -1231 4943 -1139 4949
rect -1231 4909 -1219 4943
rect -1151 4909 -1139 4943
rect -1231 4903 -1139 4909
rect -1073 4943 -981 4949
rect -1073 4909 -1061 4943
rect -993 4909 -981 4943
rect -1073 4903 -981 4909
rect -915 4943 -823 4949
rect -915 4909 -903 4943
rect -835 4909 -823 4943
rect -915 4903 -823 4909
rect -757 4943 -665 4949
rect -757 4909 -745 4943
rect -677 4909 -665 4943
rect -757 4903 -665 4909
rect -599 4943 -507 4949
rect -599 4909 -587 4943
rect -519 4909 -507 4943
rect -599 4903 -507 4909
rect -441 4943 -349 4949
rect -441 4909 -429 4943
rect -361 4909 -349 4943
rect -441 4903 -349 4909
rect -283 4943 -191 4949
rect -283 4909 -271 4943
rect -203 4909 -191 4943
rect -283 4903 -191 4909
rect -125 4943 -33 4949
rect -125 4909 -113 4943
rect -45 4909 -33 4943
rect -125 4903 -33 4909
rect 33 4943 125 4949
rect 33 4909 45 4943
rect 113 4909 125 4943
rect 33 4903 125 4909
rect 191 4943 283 4949
rect 191 4909 203 4943
rect 271 4909 283 4943
rect 191 4903 283 4909
rect 349 4943 441 4949
rect 349 4909 361 4943
rect 429 4909 441 4943
rect 349 4903 441 4909
rect 507 4943 599 4949
rect 507 4909 519 4943
rect 587 4909 599 4943
rect 507 4903 599 4909
rect 665 4943 757 4949
rect 665 4909 677 4943
rect 745 4909 757 4943
rect 665 4903 757 4909
rect 823 4943 915 4949
rect 823 4909 835 4943
rect 903 4909 915 4943
rect 823 4903 915 4909
rect 981 4943 1073 4949
rect 981 4909 993 4943
rect 1061 4909 1073 4943
rect 981 4903 1073 4909
rect 1139 4943 1231 4949
rect 1139 4909 1151 4943
rect 1219 4909 1231 4943
rect 1139 4903 1231 4909
rect 1297 4943 1389 4949
rect 1297 4909 1309 4943
rect 1377 4909 1389 4943
rect 1297 4903 1389 4909
rect 1455 4943 1547 4949
rect 1455 4909 1467 4943
rect 1535 4909 1547 4943
rect 1455 4903 1547 4909
rect -1547 4835 -1455 4841
rect -1547 4801 -1535 4835
rect -1467 4801 -1455 4835
rect -1547 4795 -1455 4801
rect -1389 4835 -1297 4841
rect -1389 4801 -1377 4835
rect -1309 4801 -1297 4835
rect -1389 4795 -1297 4801
rect -1231 4835 -1139 4841
rect -1231 4801 -1219 4835
rect -1151 4801 -1139 4835
rect -1231 4795 -1139 4801
rect -1073 4835 -981 4841
rect -1073 4801 -1061 4835
rect -993 4801 -981 4835
rect -1073 4795 -981 4801
rect -915 4835 -823 4841
rect -915 4801 -903 4835
rect -835 4801 -823 4835
rect -915 4795 -823 4801
rect -757 4835 -665 4841
rect -757 4801 -745 4835
rect -677 4801 -665 4835
rect -757 4795 -665 4801
rect -599 4835 -507 4841
rect -599 4801 -587 4835
rect -519 4801 -507 4835
rect -599 4795 -507 4801
rect -441 4835 -349 4841
rect -441 4801 -429 4835
rect -361 4801 -349 4835
rect -441 4795 -349 4801
rect -283 4835 -191 4841
rect -283 4801 -271 4835
rect -203 4801 -191 4835
rect -283 4795 -191 4801
rect -125 4835 -33 4841
rect -125 4801 -113 4835
rect -45 4801 -33 4835
rect -125 4795 -33 4801
rect 33 4835 125 4841
rect 33 4801 45 4835
rect 113 4801 125 4835
rect 33 4795 125 4801
rect 191 4835 283 4841
rect 191 4801 203 4835
rect 271 4801 283 4835
rect 191 4795 283 4801
rect 349 4835 441 4841
rect 349 4801 361 4835
rect 429 4801 441 4835
rect 349 4795 441 4801
rect 507 4835 599 4841
rect 507 4801 519 4835
rect 587 4801 599 4835
rect 507 4795 599 4801
rect 665 4835 757 4841
rect 665 4801 677 4835
rect 745 4801 757 4835
rect 665 4795 757 4801
rect 823 4835 915 4841
rect 823 4801 835 4835
rect 903 4801 915 4835
rect 823 4795 915 4801
rect 981 4835 1073 4841
rect 981 4801 993 4835
rect 1061 4801 1073 4835
rect 981 4795 1073 4801
rect 1139 4835 1231 4841
rect 1139 4801 1151 4835
rect 1219 4801 1231 4835
rect 1139 4795 1231 4801
rect 1297 4835 1389 4841
rect 1297 4801 1309 4835
rect 1377 4801 1389 4835
rect 1297 4795 1389 4801
rect 1455 4835 1547 4841
rect 1455 4801 1467 4835
rect 1535 4801 1547 4835
rect 1455 4795 1547 4801
rect -1603 4751 -1557 4763
rect -1603 3775 -1597 4751
rect -1563 3775 -1557 4751
rect -1603 3763 -1557 3775
rect -1445 4751 -1399 4763
rect -1445 3775 -1439 4751
rect -1405 3775 -1399 4751
rect -1445 3763 -1399 3775
rect -1287 4751 -1241 4763
rect -1287 3775 -1281 4751
rect -1247 3775 -1241 4751
rect -1287 3763 -1241 3775
rect -1129 4751 -1083 4763
rect -1129 3775 -1123 4751
rect -1089 3775 -1083 4751
rect -1129 3763 -1083 3775
rect -971 4751 -925 4763
rect -971 3775 -965 4751
rect -931 3775 -925 4751
rect -971 3763 -925 3775
rect -813 4751 -767 4763
rect -813 3775 -807 4751
rect -773 3775 -767 4751
rect -813 3763 -767 3775
rect -655 4751 -609 4763
rect -655 3775 -649 4751
rect -615 3775 -609 4751
rect -655 3763 -609 3775
rect -497 4751 -451 4763
rect -497 3775 -491 4751
rect -457 3775 -451 4751
rect -497 3763 -451 3775
rect -339 4751 -293 4763
rect -339 3775 -333 4751
rect -299 3775 -293 4751
rect -339 3763 -293 3775
rect -181 4751 -135 4763
rect -181 3775 -175 4751
rect -141 3775 -135 4751
rect -181 3763 -135 3775
rect -23 4751 23 4763
rect -23 3775 -17 4751
rect 17 3775 23 4751
rect -23 3763 23 3775
rect 135 4751 181 4763
rect 135 3775 141 4751
rect 175 3775 181 4751
rect 135 3763 181 3775
rect 293 4751 339 4763
rect 293 3775 299 4751
rect 333 3775 339 4751
rect 293 3763 339 3775
rect 451 4751 497 4763
rect 451 3775 457 4751
rect 491 3775 497 4751
rect 451 3763 497 3775
rect 609 4751 655 4763
rect 609 3775 615 4751
rect 649 3775 655 4751
rect 609 3763 655 3775
rect 767 4751 813 4763
rect 767 3775 773 4751
rect 807 3775 813 4751
rect 767 3763 813 3775
rect 925 4751 971 4763
rect 925 3775 931 4751
rect 965 3775 971 4751
rect 925 3763 971 3775
rect 1083 4751 1129 4763
rect 1083 3775 1089 4751
rect 1123 3775 1129 4751
rect 1083 3763 1129 3775
rect 1241 4751 1287 4763
rect 1241 3775 1247 4751
rect 1281 3775 1287 4751
rect 1241 3763 1287 3775
rect 1399 4751 1445 4763
rect 1399 3775 1405 4751
rect 1439 3775 1445 4751
rect 1399 3763 1445 3775
rect 1557 4751 1603 4763
rect 1557 3775 1563 4751
rect 1597 3775 1603 4751
rect 1557 3763 1603 3775
rect -1547 3725 -1455 3731
rect -1547 3691 -1535 3725
rect -1467 3691 -1455 3725
rect -1547 3685 -1455 3691
rect -1389 3725 -1297 3731
rect -1389 3691 -1377 3725
rect -1309 3691 -1297 3725
rect -1389 3685 -1297 3691
rect -1231 3725 -1139 3731
rect -1231 3691 -1219 3725
rect -1151 3691 -1139 3725
rect -1231 3685 -1139 3691
rect -1073 3725 -981 3731
rect -1073 3691 -1061 3725
rect -993 3691 -981 3725
rect -1073 3685 -981 3691
rect -915 3725 -823 3731
rect -915 3691 -903 3725
rect -835 3691 -823 3725
rect -915 3685 -823 3691
rect -757 3725 -665 3731
rect -757 3691 -745 3725
rect -677 3691 -665 3725
rect -757 3685 -665 3691
rect -599 3725 -507 3731
rect -599 3691 -587 3725
rect -519 3691 -507 3725
rect -599 3685 -507 3691
rect -441 3725 -349 3731
rect -441 3691 -429 3725
rect -361 3691 -349 3725
rect -441 3685 -349 3691
rect -283 3725 -191 3731
rect -283 3691 -271 3725
rect -203 3691 -191 3725
rect -283 3685 -191 3691
rect -125 3725 -33 3731
rect -125 3691 -113 3725
rect -45 3691 -33 3725
rect -125 3685 -33 3691
rect 33 3725 125 3731
rect 33 3691 45 3725
rect 113 3691 125 3725
rect 33 3685 125 3691
rect 191 3725 283 3731
rect 191 3691 203 3725
rect 271 3691 283 3725
rect 191 3685 283 3691
rect 349 3725 441 3731
rect 349 3691 361 3725
rect 429 3691 441 3725
rect 349 3685 441 3691
rect 507 3725 599 3731
rect 507 3691 519 3725
rect 587 3691 599 3725
rect 507 3685 599 3691
rect 665 3725 757 3731
rect 665 3691 677 3725
rect 745 3691 757 3725
rect 665 3685 757 3691
rect 823 3725 915 3731
rect 823 3691 835 3725
rect 903 3691 915 3725
rect 823 3685 915 3691
rect 981 3725 1073 3731
rect 981 3691 993 3725
rect 1061 3691 1073 3725
rect 981 3685 1073 3691
rect 1139 3725 1231 3731
rect 1139 3691 1151 3725
rect 1219 3691 1231 3725
rect 1139 3685 1231 3691
rect 1297 3725 1389 3731
rect 1297 3691 1309 3725
rect 1377 3691 1389 3725
rect 1297 3685 1389 3691
rect 1455 3725 1547 3731
rect 1455 3691 1467 3725
rect 1535 3691 1547 3725
rect 1455 3685 1547 3691
rect -1547 3617 -1455 3623
rect -1547 3583 -1535 3617
rect -1467 3583 -1455 3617
rect -1547 3577 -1455 3583
rect -1389 3617 -1297 3623
rect -1389 3583 -1377 3617
rect -1309 3583 -1297 3617
rect -1389 3577 -1297 3583
rect -1231 3617 -1139 3623
rect -1231 3583 -1219 3617
rect -1151 3583 -1139 3617
rect -1231 3577 -1139 3583
rect -1073 3617 -981 3623
rect -1073 3583 -1061 3617
rect -993 3583 -981 3617
rect -1073 3577 -981 3583
rect -915 3617 -823 3623
rect -915 3583 -903 3617
rect -835 3583 -823 3617
rect -915 3577 -823 3583
rect -757 3617 -665 3623
rect -757 3583 -745 3617
rect -677 3583 -665 3617
rect -757 3577 -665 3583
rect -599 3617 -507 3623
rect -599 3583 -587 3617
rect -519 3583 -507 3617
rect -599 3577 -507 3583
rect -441 3617 -349 3623
rect -441 3583 -429 3617
rect -361 3583 -349 3617
rect -441 3577 -349 3583
rect -283 3617 -191 3623
rect -283 3583 -271 3617
rect -203 3583 -191 3617
rect -283 3577 -191 3583
rect -125 3617 -33 3623
rect -125 3583 -113 3617
rect -45 3583 -33 3617
rect -125 3577 -33 3583
rect 33 3617 125 3623
rect 33 3583 45 3617
rect 113 3583 125 3617
rect 33 3577 125 3583
rect 191 3617 283 3623
rect 191 3583 203 3617
rect 271 3583 283 3617
rect 191 3577 283 3583
rect 349 3617 441 3623
rect 349 3583 361 3617
rect 429 3583 441 3617
rect 349 3577 441 3583
rect 507 3617 599 3623
rect 507 3583 519 3617
rect 587 3583 599 3617
rect 507 3577 599 3583
rect 665 3617 757 3623
rect 665 3583 677 3617
rect 745 3583 757 3617
rect 665 3577 757 3583
rect 823 3617 915 3623
rect 823 3583 835 3617
rect 903 3583 915 3617
rect 823 3577 915 3583
rect 981 3617 1073 3623
rect 981 3583 993 3617
rect 1061 3583 1073 3617
rect 981 3577 1073 3583
rect 1139 3617 1231 3623
rect 1139 3583 1151 3617
rect 1219 3583 1231 3617
rect 1139 3577 1231 3583
rect 1297 3617 1389 3623
rect 1297 3583 1309 3617
rect 1377 3583 1389 3617
rect 1297 3577 1389 3583
rect 1455 3617 1547 3623
rect 1455 3583 1467 3617
rect 1535 3583 1547 3617
rect 1455 3577 1547 3583
rect -1603 3533 -1557 3545
rect -1603 2557 -1597 3533
rect -1563 2557 -1557 3533
rect -1603 2545 -1557 2557
rect -1445 3533 -1399 3545
rect -1445 2557 -1439 3533
rect -1405 2557 -1399 3533
rect -1445 2545 -1399 2557
rect -1287 3533 -1241 3545
rect -1287 2557 -1281 3533
rect -1247 2557 -1241 3533
rect -1287 2545 -1241 2557
rect -1129 3533 -1083 3545
rect -1129 2557 -1123 3533
rect -1089 2557 -1083 3533
rect -1129 2545 -1083 2557
rect -971 3533 -925 3545
rect -971 2557 -965 3533
rect -931 2557 -925 3533
rect -971 2545 -925 2557
rect -813 3533 -767 3545
rect -813 2557 -807 3533
rect -773 2557 -767 3533
rect -813 2545 -767 2557
rect -655 3533 -609 3545
rect -655 2557 -649 3533
rect -615 2557 -609 3533
rect -655 2545 -609 2557
rect -497 3533 -451 3545
rect -497 2557 -491 3533
rect -457 2557 -451 3533
rect -497 2545 -451 2557
rect -339 3533 -293 3545
rect -339 2557 -333 3533
rect -299 2557 -293 3533
rect -339 2545 -293 2557
rect -181 3533 -135 3545
rect -181 2557 -175 3533
rect -141 2557 -135 3533
rect -181 2545 -135 2557
rect -23 3533 23 3545
rect -23 2557 -17 3533
rect 17 2557 23 3533
rect -23 2545 23 2557
rect 135 3533 181 3545
rect 135 2557 141 3533
rect 175 2557 181 3533
rect 135 2545 181 2557
rect 293 3533 339 3545
rect 293 2557 299 3533
rect 333 2557 339 3533
rect 293 2545 339 2557
rect 451 3533 497 3545
rect 451 2557 457 3533
rect 491 2557 497 3533
rect 451 2545 497 2557
rect 609 3533 655 3545
rect 609 2557 615 3533
rect 649 2557 655 3533
rect 609 2545 655 2557
rect 767 3533 813 3545
rect 767 2557 773 3533
rect 807 2557 813 3533
rect 767 2545 813 2557
rect 925 3533 971 3545
rect 925 2557 931 3533
rect 965 2557 971 3533
rect 925 2545 971 2557
rect 1083 3533 1129 3545
rect 1083 2557 1089 3533
rect 1123 2557 1129 3533
rect 1083 2545 1129 2557
rect 1241 3533 1287 3545
rect 1241 2557 1247 3533
rect 1281 2557 1287 3533
rect 1241 2545 1287 2557
rect 1399 3533 1445 3545
rect 1399 2557 1405 3533
rect 1439 2557 1445 3533
rect 1399 2545 1445 2557
rect 1557 3533 1603 3545
rect 1557 2557 1563 3533
rect 1597 2557 1603 3533
rect 1557 2545 1603 2557
rect -1547 2507 -1455 2513
rect -1547 2473 -1535 2507
rect -1467 2473 -1455 2507
rect -1547 2467 -1455 2473
rect -1389 2507 -1297 2513
rect -1389 2473 -1377 2507
rect -1309 2473 -1297 2507
rect -1389 2467 -1297 2473
rect -1231 2507 -1139 2513
rect -1231 2473 -1219 2507
rect -1151 2473 -1139 2507
rect -1231 2467 -1139 2473
rect -1073 2507 -981 2513
rect -1073 2473 -1061 2507
rect -993 2473 -981 2507
rect -1073 2467 -981 2473
rect -915 2507 -823 2513
rect -915 2473 -903 2507
rect -835 2473 -823 2507
rect -915 2467 -823 2473
rect -757 2507 -665 2513
rect -757 2473 -745 2507
rect -677 2473 -665 2507
rect -757 2467 -665 2473
rect -599 2507 -507 2513
rect -599 2473 -587 2507
rect -519 2473 -507 2507
rect -599 2467 -507 2473
rect -441 2507 -349 2513
rect -441 2473 -429 2507
rect -361 2473 -349 2507
rect -441 2467 -349 2473
rect -283 2507 -191 2513
rect -283 2473 -271 2507
rect -203 2473 -191 2507
rect -283 2467 -191 2473
rect -125 2507 -33 2513
rect -125 2473 -113 2507
rect -45 2473 -33 2507
rect -125 2467 -33 2473
rect 33 2507 125 2513
rect 33 2473 45 2507
rect 113 2473 125 2507
rect 33 2467 125 2473
rect 191 2507 283 2513
rect 191 2473 203 2507
rect 271 2473 283 2507
rect 191 2467 283 2473
rect 349 2507 441 2513
rect 349 2473 361 2507
rect 429 2473 441 2507
rect 349 2467 441 2473
rect 507 2507 599 2513
rect 507 2473 519 2507
rect 587 2473 599 2507
rect 507 2467 599 2473
rect 665 2507 757 2513
rect 665 2473 677 2507
rect 745 2473 757 2507
rect 665 2467 757 2473
rect 823 2507 915 2513
rect 823 2473 835 2507
rect 903 2473 915 2507
rect 823 2467 915 2473
rect 981 2507 1073 2513
rect 981 2473 993 2507
rect 1061 2473 1073 2507
rect 981 2467 1073 2473
rect 1139 2507 1231 2513
rect 1139 2473 1151 2507
rect 1219 2473 1231 2507
rect 1139 2467 1231 2473
rect 1297 2507 1389 2513
rect 1297 2473 1309 2507
rect 1377 2473 1389 2507
rect 1297 2467 1389 2473
rect 1455 2507 1547 2513
rect 1455 2473 1467 2507
rect 1535 2473 1547 2507
rect 1455 2467 1547 2473
rect -1547 2399 -1455 2405
rect -1547 2365 -1535 2399
rect -1467 2365 -1455 2399
rect -1547 2359 -1455 2365
rect -1389 2399 -1297 2405
rect -1389 2365 -1377 2399
rect -1309 2365 -1297 2399
rect -1389 2359 -1297 2365
rect -1231 2399 -1139 2405
rect -1231 2365 -1219 2399
rect -1151 2365 -1139 2399
rect -1231 2359 -1139 2365
rect -1073 2399 -981 2405
rect -1073 2365 -1061 2399
rect -993 2365 -981 2399
rect -1073 2359 -981 2365
rect -915 2399 -823 2405
rect -915 2365 -903 2399
rect -835 2365 -823 2399
rect -915 2359 -823 2365
rect -757 2399 -665 2405
rect -757 2365 -745 2399
rect -677 2365 -665 2399
rect -757 2359 -665 2365
rect -599 2399 -507 2405
rect -599 2365 -587 2399
rect -519 2365 -507 2399
rect -599 2359 -507 2365
rect -441 2399 -349 2405
rect -441 2365 -429 2399
rect -361 2365 -349 2399
rect -441 2359 -349 2365
rect -283 2399 -191 2405
rect -283 2365 -271 2399
rect -203 2365 -191 2399
rect -283 2359 -191 2365
rect -125 2399 -33 2405
rect -125 2365 -113 2399
rect -45 2365 -33 2399
rect -125 2359 -33 2365
rect 33 2399 125 2405
rect 33 2365 45 2399
rect 113 2365 125 2399
rect 33 2359 125 2365
rect 191 2399 283 2405
rect 191 2365 203 2399
rect 271 2365 283 2399
rect 191 2359 283 2365
rect 349 2399 441 2405
rect 349 2365 361 2399
rect 429 2365 441 2399
rect 349 2359 441 2365
rect 507 2399 599 2405
rect 507 2365 519 2399
rect 587 2365 599 2399
rect 507 2359 599 2365
rect 665 2399 757 2405
rect 665 2365 677 2399
rect 745 2365 757 2399
rect 665 2359 757 2365
rect 823 2399 915 2405
rect 823 2365 835 2399
rect 903 2365 915 2399
rect 823 2359 915 2365
rect 981 2399 1073 2405
rect 981 2365 993 2399
rect 1061 2365 1073 2399
rect 981 2359 1073 2365
rect 1139 2399 1231 2405
rect 1139 2365 1151 2399
rect 1219 2365 1231 2399
rect 1139 2359 1231 2365
rect 1297 2399 1389 2405
rect 1297 2365 1309 2399
rect 1377 2365 1389 2399
rect 1297 2359 1389 2365
rect 1455 2399 1547 2405
rect 1455 2365 1467 2399
rect 1535 2365 1547 2399
rect 1455 2359 1547 2365
rect -1603 2315 -1557 2327
rect -1603 1339 -1597 2315
rect -1563 1339 -1557 2315
rect -1603 1327 -1557 1339
rect -1445 2315 -1399 2327
rect -1445 1339 -1439 2315
rect -1405 1339 -1399 2315
rect -1445 1327 -1399 1339
rect -1287 2315 -1241 2327
rect -1287 1339 -1281 2315
rect -1247 1339 -1241 2315
rect -1287 1327 -1241 1339
rect -1129 2315 -1083 2327
rect -1129 1339 -1123 2315
rect -1089 1339 -1083 2315
rect -1129 1327 -1083 1339
rect -971 2315 -925 2327
rect -971 1339 -965 2315
rect -931 1339 -925 2315
rect -971 1327 -925 1339
rect -813 2315 -767 2327
rect -813 1339 -807 2315
rect -773 1339 -767 2315
rect -813 1327 -767 1339
rect -655 2315 -609 2327
rect -655 1339 -649 2315
rect -615 1339 -609 2315
rect -655 1327 -609 1339
rect -497 2315 -451 2327
rect -497 1339 -491 2315
rect -457 1339 -451 2315
rect -497 1327 -451 1339
rect -339 2315 -293 2327
rect -339 1339 -333 2315
rect -299 1339 -293 2315
rect -339 1327 -293 1339
rect -181 2315 -135 2327
rect -181 1339 -175 2315
rect -141 1339 -135 2315
rect -181 1327 -135 1339
rect -23 2315 23 2327
rect -23 1339 -17 2315
rect 17 1339 23 2315
rect -23 1327 23 1339
rect 135 2315 181 2327
rect 135 1339 141 2315
rect 175 1339 181 2315
rect 135 1327 181 1339
rect 293 2315 339 2327
rect 293 1339 299 2315
rect 333 1339 339 2315
rect 293 1327 339 1339
rect 451 2315 497 2327
rect 451 1339 457 2315
rect 491 1339 497 2315
rect 451 1327 497 1339
rect 609 2315 655 2327
rect 609 1339 615 2315
rect 649 1339 655 2315
rect 609 1327 655 1339
rect 767 2315 813 2327
rect 767 1339 773 2315
rect 807 1339 813 2315
rect 767 1327 813 1339
rect 925 2315 971 2327
rect 925 1339 931 2315
rect 965 1339 971 2315
rect 925 1327 971 1339
rect 1083 2315 1129 2327
rect 1083 1339 1089 2315
rect 1123 1339 1129 2315
rect 1083 1327 1129 1339
rect 1241 2315 1287 2327
rect 1241 1339 1247 2315
rect 1281 1339 1287 2315
rect 1241 1327 1287 1339
rect 1399 2315 1445 2327
rect 1399 1339 1405 2315
rect 1439 1339 1445 2315
rect 1399 1327 1445 1339
rect 1557 2315 1603 2327
rect 1557 1339 1563 2315
rect 1597 1339 1603 2315
rect 1557 1327 1603 1339
rect -1547 1289 -1455 1295
rect -1547 1255 -1535 1289
rect -1467 1255 -1455 1289
rect -1547 1249 -1455 1255
rect -1389 1289 -1297 1295
rect -1389 1255 -1377 1289
rect -1309 1255 -1297 1289
rect -1389 1249 -1297 1255
rect -1231 1289 -1139 1295
rect -1231 1255 -1219 1289
rect -1151 1255 -1139 1289
rect -1231 1249 -1139 1255
rect -1073 1289 -981 1295
rect -1073 1255 -1061 1289
rect -993 1255 -981 1289
rect -1073 1249 -981 1255
rect -915 1289 -823 1295
rect -915 1255 -903 1289
rect -835 1255 -823 1289
rect -915 1249 -823 1255
rect -757 1289 -665 1295
rect -757 1255 -745 1289
rect -677 1255 -665 1289
rect -757 1249 -665 1255
rect -599 1289 -507 1295
rect -599 1255 -587 1289
rect -519 1255 -507 1289
rect -599 1249 -507 1255
rect -441 1289 -349 1295
rect -441 1255 -429 1289
rect -361 1255 -349 1289
rect -441 1249 -349 1255
rect -283 1289 -191 1295
rect -283 1255 -271 1289
rect -203 1255 -191 1289
rect -283 1249 -191 1255
rect -125 1289 -33 1295
rect -125 1255 -113 1289
rect -45 1255 -33 1289
rect -125 1249 -33 1255
rect 33 1289 125 1295
rect 33 1255 45 1289
rect 113 1255 125 1289
rect 33 1249 125 1255
rect 191 1289 283 1295
rect 191 1255 203 1289
rect 271 1255 283 1289
rect 191 1249 283 1255
rect 349 1289 441 1295
rect 349 1255 361 1289
rect 429 1255 441 1289
rect 349 1249 441 1255
rect 507 1289 599 1295
rect 507 1255 519 1289
rect 587 1255 599 1289
rect 507 1249 599 1255
rect 665 1289 757 1295
rect 665 1255 677 1289
rect 745 1255 757 1289
rect 665 1249 757 1255
rect 823 1289 915 1295
rect 823 1255 835 1289
rect 903 1255 915 1289
rect 823 1249 915 1255
rect 981 1289 1073 1295
rect 981 1255 993 1289
rect 1061 1255 1073 1289
rect 981 1249 1073 1255
rect 1139 1289 1231 1295
rect 1139 1255 1151 1289
rect 1219 1255 1231 1289
rect 1139 1249 1231 1255
rect 1297 1289 1389 1295
rect 1297 1255 1309 1289
rect 1377 1255 1389 1289
rect 1297 1249 1389 1255
rect 1455 1289 1547 1295
rect 1455 1255 1467 1289
rect 1535 1255 1547 1289
rect 1455 1249 1547 1255
rect -1547 1181 -1455 1187
rect -1547 1147 -1535 1181
rect -1467 1147 -1455 1181
rect -1547 1141 -1455 1147
rect -1389 1181 -1297 1187
rect -1389 1147 -1377 1181
rect -1309 1147 -1297 1181
rect -1389 1141 -1297 1147
rect -1231 1181 -1139 1187
rect -1231 1147 -1219 1181
rect -1151 1147 -1139 1181
rect -1231 1141 -1139 1147
rect -1073 1181 -981 1187
rect -1073 1147 -1061 1181
rect -993 1147 -981 1181
rect -1073 1141 -981 1147
rect -915 1181 -823 1187
rect -915 1147 -903 1181
rect -835 1147 -823 1181
rect -915 1141 -823 1147
rect -757 1181 -665 1187
rect -757 1147 -745 1181
rect -677 1147 -665 1181
rect -757 1141 -665 1147
rect -599 1181 -507 1187
rect -599 1147 -587 1181
rect -519 1147 -507 1181
rect -599 1141 -507 1147
rect -441 1181 -349 1187
rect -441 1147 -429 1181
rect -361 1147 -349 1181
rect -441 1141 -349 1147
rect -283 1181 -191 1187
rect -283 1147 -271 1181
rect -203 1147 -191 1181
rect -283 1141 -191 1147
rect -125 1181 -33 1187
rect -125 1147 -113 1181
rect -45 1147 -33 1181
rect -125 1141 -33 1147
rect 33 1181 125 1187
rect 33 1147 45 1181
rect 113 1147 125 1181
rect 33 1141 125 1147
rect 191 1181 283 1187
rect 191 1147 203 1181
rect 271 1147 283 1181
rect 191 1141 283 1147
rect 349 1181 441 1187
rect 349 1147 361 1181
rect 429 1147 441 1181
rect 349 1141 441 1147
rect 507 1181 599 1187
rect 507 1147 519 1181
rect 587 1147 599 1181
rect 507 1141 599 1147
rect 665 1181 757 1187
rect 665 1147 677 1181
rect 745 1147 757 1181
rect 665 1141 757 1147
rect 823 1181 915 1187
rect 823 1147 835 1181
rect 903 1147 915 1181
rect 823 1141 915 1147
rect 981 1181 1073 1187
rect 981 1147 993 1181
rect 1061 1147 1073 1181
rect 981 1141 1073 1147
rect 1139 1181 1231 1187
rect 1139 1147 1151 1181
rect 1219 1147 1231 1181
rect 1139 1141 1231 1147
rect 1297 1181 1389 1187
rect 1297 1147 1309 1181
rect 1377 1147 1389 1181
rect 1297 1141 1389 1147
rect 1455 1181 1547 1187
rect 1455 1147 1467 1181
rect 1535 1147 1547 1181
rect 1455 1141 1547 1147
rect -1603 1097 -1557 1109
rect -1603 121 -1597 1097
rect -1563 121 -1557 1097
rect -1603 109 -1557 121
rect -1445 1097 -1399 1109
rect -1445 121 -1439 1097
rect -1405 121 -1399 1097
rect -1445 109 -1399 121
rect -1287 1097 -1241 1109
rect -1287 121 -1281 1097
rect -1247 121 -1241 1097
rect -1287 109 -1241 121
rect -1129 1097 -1083 1109
rect -1129 121 -1123 1097
rect -1089 121 -1083 1097
rect -1129 109 -1083 121
rect -971 1097 -925 1109
rect -971 121 -965 1097
rect -931 121 -925 1097
rect -971 109 -925 121
rect -813 1097 -767 1109
rect -813 121 -807 1097
rect -773 121 -767 1097
rect -813 109 -767 121
rect -655 1097 -609 1109
rect -655 121 -649 1097
rect -615 121 -609 1097
rect -655 109 -609 121
rect -497 1097 -451 1109
rect -497 121 -491 1097
rect -457 121 -451 1097
rect -497 109 -451 121
rect -339 1097 -293 1109
rect -339 121 -333 1097
rect -299 121 -293 1097
rect -339 109 -293 121
rect -181 1097 -135 1109
rect -181 121 -175 1097
rect -141 121 -135 1097
rect -181 109 -135 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 135 1097 181 1109
rect 135 121 141 1097
rect 175 121 181 1097
rect 135 109 181 121
rect 293 1097 339 1109
rect 293 121 299 1097
rect 333 121 339 1097
rect 293 109 339 121
rect 451 1097 497 1109
rect 451 121 457 1097
rect 491 121 497 1097
rect 451 109 497 121
rect 609 1097 655 1109
rect 609 121 615 1097
rect 649 121 655 1097
rect 609 109 655 121
rect 767 1097 813 1109
rect 767 121 773 1097
rect 807 121 813 1097
rect 767 109 813 121
rect 925 1097 971 1109
rect 925 121 931 1097
rect 965 121 971 1097
rect 925 109 971 121
rect 1083 1097 1129 1109
rect 1083 121 1089 1097
rect 1123 121 1129 1097
rect 1083 109 1129 121
rect 1241 1097 1287 1109
rect 1241 121 1247 1097
rect 1281 121 1287 1097
rect 1241 109 1287 121
rect 1399 1097 1445 1109
rect 1399 121 1405 1097
rect 1439 121 1445 1097
rect 1399 109 1445 121
rect 1557 1097 1603 1109
rect 1557 121 1563 1097
rect 1597 121 1603 1097
rect 1557 109 1603 121
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect -1603 -121 -1557 -109
rect -1603 -1097 -1597 -121
rect -1563 -1097 -1557 -121
rect -1603 -1109 -1557 -1097
rect -1445 -121 -1399 -109
rect -1445 -1097 -1439 -121
rect -1405 -1097 -1399 -121
rect -1445 -1109 -1399 -1097
rect -1287 -121 -1241 -109
rect -1287 -1097 -1281 -121
rect -1247 -1097 -1241 -121
rect -1287 -1109 -1241 -1097
rect -1129 -121 -1083 -109
rect -1129 -1097 -1123 -121
rect -1089 -1097 -1083 -121
rect -1129 -1109 -1083 -1097
rect -971 -121 -925 -109
rect -971 -1097 -965 -121
rect -931 -1097 -925 -121
rect -971 -1109 -925 -1097
rect -813 -121 -767 -109
rect -813 -1097 -807 -121
rect -773 -1097 -767 -121
rect -813 -1109 -767 -1097
rect -655 -121 -609 -109
rect -655 -1097 -649 -121
rect -615 -1097 -609 -121
rect -655 -1109 -609 -1097
rect -497 -121 -451 -109
rect -497 -1097 -491 -121
rect -457 -1097 -451 -121
rect -497 -1109 -451 -1097
rect -339 -121 -293 -109
rect -339 -1097 -333 -121
rect -299 -1097 -293 -121
rect -339 -1109 -293 -1097
rect -181 -121 -135 -109
rect -181 -1097 -175 -121
rect -141 -1097 -135 -121
rect -181 -1109 -135 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 135 -121 181 -109
rect 135 -1097 141 -121
rect 175 -1097 181 -121
rect 135 -1109 181 -1097
rect 293 -121 339 -109
rect 293 -1097 299 -121
rect 333 -1097 339 -121
rect 293 -1109 339 -1097
rect 451 -121 497 -109
rect 451 -1097 457 -121
rect 491 -1097 497 -121
rect 451 -1109 497 -1097
rect 609 -121 655 -109
rect 609 -1097 615 -121
rect 649 -1097 655 -121
rect 609 -1109 655 -1097
rect 767 -121 813 -109
rect 767 -1097 773 -121
rect 807 -1097 813 -121
rect 767 -1109 813 -1097
rect 925 -121 971 -109
rect 925 -1097 931 -121
rect 965 -1097 971 -121
rect 925 -1109 971 -1097
rect 1083 -121 1129 -109
rect 1083 -1097 1089 -121
rect 1123 -1097 1129 -121
rect 1083 -1109 1129 -1097
rect 1241 -121 1287 -109
rect 1241 -1097 1247 -121
rect 1281 -1097 1287 -121
rect 1241 -1109 1287 -1097
rect 1399 -121 1445 -109
rect 1399 -1097 1405 -121
rect 1439 -1097 1445 -121
rect 1399 -1109 1445 -1097
rect 1557 -121 1603 -109
rect 1557 -1097 1563 -121
rect 1597 -1097 1603 -121
rect 1557 -1109 1603 -1097
rect -1547 -1147 -1455 -1141
rect -1547 -1181 -1535 -1147
rect -1467 -1181 -1455 -1147
rect -1547 -1187 -1455 -1181
rect -1389 -1147 -1297 -1141
rect -1389 -1181 -1377 -1147
rect -1309 -1181 -1297 -1147
rect -1389 -1187 -1297 -1181
rect -1231 -1147 -1139 -1141
rect -1231 -1181 -1219 -1147
rect -1151 -1181 -1139 -1147
rect -1231 -1187 -1139 -1181
rect -1073 -1147 -981 -1141
rect -1073 -1181 -1061 -1147
rect -993 -1181 -981 -1147
rect -1073 -1187 -981 -1181
rect -915 -1147 -823 -1141
rect -915 -1181 -903 -1147
rect -835 -1181 -823 -1147
rect -915 -1187 -823 -1181
rect -757 -1147 -665 -1141
rect -757 -1181 -745 -1147
rect -677 -1181 -665 -1147
rect -757 -1187 -665 -1181
rect -599 -1147 -507 -1141
rect -599 -1181 -587 -1147
rect -519 -1181 -507 -1147
rect -599 -1187 -507 -1181
rect -441 -1147 -349 -1141
rect -441 -1181 -429 -1147
rect -361 -1181 -349 -1147
rect -441 -1187 -349 -1181
rect -283 -1147 -191 -1141
rect -283 -1181 -271 -1147
rect -203 -1181 -191 -1147
rect -283 -1187 -191 -1181
rect -125 -1147 -33 -1141
rect -125 -1181 -113 -1147
rect -45 -1181 -33 -1147
rect -125 -1187 -33 -1181
rect 33 -1147 125 -1141
rect 33 -1181 45 -1147
rect 113 -1181 125 -1147
rect 33 -1187 125 -1181
rect 191 -1147 283 -1141
rect 191 -1181 203 -1147
rect 271 -1181 283 -1147
rect 191 -1187 283 -1181
rect 349 -1147 441 -1141
rect 349 -1181 361 -1147
rect 429 -1181 441 -1147
rect 349 -1187 441 -1181
rect 507 -1147 599 -1141
rect 507 -1181 519 -1147
rect 587 -1181 599 -1147
rect 507 -1187 599 -1181
rect 665 -1147 757 -1141
rect 665 -1181 677 -1147
rect 745 -1181 757 -1147
rect 665 -1187 757 -1181
rect 823 -1147 915 -1141
rect 823 -1181 835 -1147
rect 903 -1181 915 -1147
rect 823 -1187 915 -1181
rect 981 -1147 1073 -1141
rect 981 -1181 993 -1147
rect 1061 -1181 1073 -1147
rect 981 -1187 1073 -1181
rect 1139 -1147 1231 -1141
rect 1139 -1181 1151 -1147
rect 1219 -1181 1231 -1147
rect 1139 -1187 1231 -1181
rect 1297 -1147 1389 -1141
rect 1297 -1181 1309 -1147
rect 1377 -1181 1389 -1147
rect 1297 -1187 1389 -1181
rect 1455 -1147 1547 -1141
rect 1455 -1181 1467 -1147
rect 1535 -1181 1547 -1147
rect 1455 -1187 1547 -1181
rect -1547 -1255 -1455 -1249
rect -1547 -1289 -1535 -1255
rect -1467 -1289 -1455 -1255
rect -1547 -1295 -1455 -1289
rect -1389 -1255 -1297 -1249
rect -1389 -1289 -1377 -1255
rect -1309 -1289 -1297 -1255
rect -1389 -1295 -1297 -1289
rect -1231 -1255 -1139 -1249
rect -1231 -1289 -1219 -1255
rect -1151 -1289 -1139 -1255
rect -1231 -1295 -1139 -1289
rect -1073 -1255 -981 -1249
rect -1073 -1289 -1061 -1255
rect -993 -1289 -981 -1255
rect -1073 -1295 -981 -1289
rect -915 -1255 -823 -1249
rect -915 -1289 -903 -1255
rect -835 -1289 -823 -1255
rect -915 -1295 -823 -1289
rect -757 -1255 -665 -1249
rect -757 -1289 -745 -1255
rect -677 -1289 -665 -1255
rect -757 -1295 -665 -1289
rect -599 -1255 -507 -1249
rect -599 -1289 -587 -1255
rect -519 -1289 -507 -1255
rect -599 -1295 -507 -1289
rect -441 -1255 -349 -1249
rect -441 -1289 -429 -1255
rect -361 -1289 -349 -1255
rect -441 -1295 -349 -1289
rect -283 -1255 -191 -1249
rect -283 -1289 -271 -1255
rect -203 -1289 -191 -1255
rect -283 -1295 -191 -1289
rect -125 -1255 -33 -1249
rect -125 -1289 -113 -1255
rect -45 -1289 -33 -1255
rect -125 -1295 -33 -1289
rect 33 -1255 125 -1249
rect 33 -1289 45 -1255
rect 113 -1289 125 -1255
rect 33 -1295 125 -1289
rect 191 -1255 283 -1249
rect 191 -1289 203 -1255
rect 271 -1289 283 -1255
rect 191 -1295 283 -1289
rect 349 -1255 441 -1249
rect 349 -1289 361 -1255
rect 429 -1289 441 -1255
rect 349 -1295 441 -1289
rect 507 -1255 599 -1249
rect 507 -1289 519 -1255
rect 587 -1289 599 -1255
rect 507 -1295 599 -1289
rect 665 -1255 757 -1249
rect 665 -1289 677 -1255
rect 745 -1289 757 -1255
rect 665 -1295 757 -1289
rect 823 -1255 915 -1249
rect 823 -1289 835 -1255
rect 903 -1289 915 -1255
rect 823 -1295 915 -1289
rect 981 -1255 1073 -1249
rect 981 -1289 993 -1255
rect 1061 -1289 1073 -1255
rect 981 -1295 1073 -1289
rect 1139 -1255 1231 -1249
rect 1139 -1289 1151 -1255
rect 1219 -1289 1231 -1255
rect 1139 -1295 1231 -1289
rect 1297 -1255 1389 -1249
rect 1297 -1289 1309 -1255
rect 1377 -1289 1389 -1255
rect 1297 -1295 1389 -1289
rect 1455 -1255 1547 -1249
rect 1455 -1289 1467 -1255
rect 1535 -1289 1547 -1255
rect 1455 -1295 1547 -1289
rect -1603 -1339 -1557 -1327
rect -1603 -2315 -1597 -1339
rect -1563 -2315 -1557 -1339
rect -1603 -2327 -1557 -2315
rect -1445 -1339 -1399 -1327
rect -1445 -2315 -1439 -1339
rect -1405 -2315 -1399 -1339
rect -1445 -2327 -1399 -2315
rect -1287 -1339 -1241 -1327
rect -1287 -2315 -1281 -1339
rect -1247 -2315 -1241 -1339
rect -1287 -2327 -1241 -2315
rect -1129 -1339 -1083 -1327
rect -1129 -2315 -1123 -1339
rect -1089 -2315 -1083 -1339
rect -1129 -2327 -1083 -2315
rect -971 -1339 -925 -1327
rect -971 -2315 -965 -1339
rect -931 -2315 -925 -1339
rect -971 -2327 -925 -2315
rect -813 -1339 -767 -1327
rect -813 -2315 -807 -1339
rect -773 -2315 -767 -1339
rect -813 -2327 -767 -2315
rect -655 -1339 -609 -1327
rect -655 -2315 -649 -1339
rect -615 -2315 -609 -1339
rect -655 -2327 -609 -2315
rect -497 -1339 -451 -1327
rect -497 -2315 -491 -1339
rect -457 -2315 -451 -1339
rect -497 -2327 -451 -2315
rect -339 -1339 -293 -1327
rect -339 -2315 -333 -1339
rect -299 -2315 -293 -1339
rect -339 -2327 -293 -2315
rect -181 -1339 -135 -1327
rect -181 -2315 -175 -1339
rect -141 -2315 -135 -1339
rect -181 -2327 -135 -2315
rect -23 -1339 23 -1327
rect -23 -2315 -17 -1339
rect 17 -2315 23 -1339
rect -23 -2327 23 -2315
rect 135 -1339 181 -1327
rect 135 -2315 141 -1339
rect 175 -2315 181 -1339
rect 135 -2327 181 -2315
rect 293 -1339 339 -1327
rect 293 -2315 299 -1339
rect 333 -2315 339 -1339
rect 293 -2327 339 -2315
rect 451 -1339 497 -1327
rect 451 -2315 457 -1339
rect 491 -2315 497 -1339
rect 451 -2327 497 -2315
rect 609 -1339 655 -1327
rect 609 -2315 615 -1339
rect 649 -2315 655 -1339
rect 609 -2327 655 -2315
rect 767 -1339 813 -1327
rect 767 -2315 773 -1339
rect 807 -2315 813 -1339
rect 767 -2327 813 -2315
rect 925 -1339 971 -1327
rect 925 -2315 931 -1339
rect 965 -2315 971 -1339
rect 925 -2327 971 -2315
rect 1083 -1339 1129 -1327
rect 1083 -2315 1089 -1339
rect 1123 -2315 1129 -1339
rect 1083 -2327 1129 -2315
rect 1241 -1339 1287 -1327
rect 1241 -2315 1247 -1339
rect 1281 -2315 1287 -1339
rect 1241 -2327 1287 -2315
rect 1399 -1339 1445 -1327
rect 1399 -2315 1405 -1339
rect 1439 -2315 1445 -1339
rect 1399 -2327 1445 -2315
rect 1557 -1339 1603 -1327
rect 1557 -2315 1563 -1339
rect 1597 -2315 1603 -1339
rect 1557 -2327 1603 -2315
rect -1547 -2365 -1455 -2359
rect -1547 -2399 -1535 -2365
rect -1467 -2399 -1455 -2365
rect -1547 -2405 -1455 -2399
rect -1389 -2365 -1297 -2359
rect -1389 -2399 -1377 -2365
rect -1309 -2399 -1297 -2365
rect -1389 -2405 -1297 -2399
rect -1231 -2365 -1139 -2359
rect -1231 -2399 -1219 -2365
rect -1151 -2399 -1139 -2365
rect -1231 -2405 -1139 -2399
rect -1073 -2365 -981 -2359
rect -1073 -2399 -1061 -2365
rect -993 -2399 -981 -2365
rect -1073 -2405 -981 -2399
rect -915 -2365 -823 -2359
rect -915 -2399 -903 -2365
rect -835 -2399 -823 -2365
rect -915 -2405 -823 -2399
rect -757 -2365 -665 -2359
rect -757 -2399 -745 -2365
rect -677 -2399 -665 -2365
rect -757 -2405 -665 -2399
rect -599 -2365 -507 -2359
rect -599 -2399 -587 -2365
rect -519 -2399 -507 -2365
rect -599 -2405 -507 -2399
rect -441 -2365 -349 -2359
rect -441 -2399 -429 -2365
rect -361 -2399 -349 -2365
rect -441 -2405 -349 -2399
rect -283 -2365 -191 -2359
rect -283 -2399 -271 -2365
rect -203 -2399 -191 -2365
rect -283 -2405 -191 -2399
rect -125 -2365 -33 -2359
rect -125 -2399 -113 -2365
rect -45 -2399 -33 -2365
rect -125 -2405 -33 -2399
rect 33 -2365 125 -2359
rect 33 -2399 45 -2365
rect 113 -2399 125 -2365
rect 33 -2405 125 -2399
rect 191 -2365 283 -2359
rect 191 -2399 203 -2365
rect 271 -2399 283 -2365
rect 191 -2405 283 -2399
rect 349 -2365 441 -2359
rect 349 -2399 361 -2365
rect 429 -2399 441 -2365
rect 349 -2405 441 -2399
rect 507 -2365 599 -2359
rect 507 -2399 519 -2365
rect 587 -2399 599 -2365
rect 507 -2405 599 -2399
rect 665 -2365 757 -2359
rect 665 -2399 677 -2365
rect 745 -2399 757 -2365
rect 665 -2405 757 -2399
rect 823 -2365 915 -2359
rect 823 -2399 835 -2365
rect 903 -2399 915 -2365
rect 823 -2405 915 -2399
rect 981 -2365 1073 -2359
rect 981 -2399 993 -2365
rect 1061 -2399 1073 -2365
rect 981 -2405 1073 -2399
rect 1139 -2365 1231 -2359
rect 1139 -2399 1151 -2365
rect 1219 -2399 1231 -2365
rect 1139 -2405 1231 -2399
rect 1297 -2365 1389 -2359
rect 1297 -2399 1309 -2365
rect 1377 -2399 1389 -2365
rect 1297 -2405 1389 -2399
rect 1455 -2365 1547 -2359
rect 1455 -2399 1467 -2365
rect 1535 -2399 1547 -2365
rect 1455 -2405 1547 -2399
rect -1547 -2473 -1455 -2467
rect -1547 -2507 -1535 -2473
rect -1467 -2507 -1455 -2473
rect -1547 -2513 -1455 -2507
rect -1389 -2473 -1297 -2467
rect -1389 -2507 -1377 -2473
rect -1309 -2507 -1297 -2473
rect -1389 -2513 -1297 -2507
rect -1231 -2473 -1139 -2467
rect -1231 -2507 -1219 -2473
rect -1151 -2507 -1139 -2473
rect -1231 -2513 -1139 -2507
rect -1073 -2473 -981 -2467
rect -1073 -2507 -1061 -2473
rect -993 -2507 -981 -2473
rect -1073 -2513 -981 -2507
rect -915 -2473 -823 -2467
rect -915 -2507 -903 -2473
rect -835 -2507 -823 -2473
rect -915 -2513 -823 -2507
rect -757 -2473 -665 -2467
rect -757 -2507 -745 -2473
rect -677 -2507 -665 -2473
rect -757 -2513 -665 -2507
rect -599 -2473 -507 -2467
rect -599 -2507 -587 -2473
rect -519 -2507 -507 -2473
rect -599 -2513 -507 -2507
rect -441 -2473 -349 -2467
rect -441 -2507 -429 -2473
rect -361 -2507 -349 -2473
rect -441 -2513 -349 -2507
rect -283 -2473 -191 -2467
rect -283 -2507 -271 -2473
rect -203 -2507 -191 -2473
rect -283 -2513 -191 -2507
rect -125 -2473 -33 -2467
rect -125 -2507 -113 -2473
rect -45 -2507 -33 -2473
rect -125 -2513 -33 -2507
rect 33 -2473 125 -2467
rect 33 -2507 45 -2473
rect 113 -2507 125 -2473
rect 33 -2513 125 -2507
rect 191 -2473 283 -2467
rect 191 -2507 203 -2473
rect 271 -2507 283 -2473
rect 191 -2513 283 -2507
rect 349 -2473 441 -2467
rect 349 -2507 361 -2473
rect 429 -2507 441 -2473
rect 349 -2513 441 -2507
rect 507 -2473 599 -2467
rect 507 -2507 519 -2473
rect 587 -2507 599 -2473
rect 507 -2513 599 -2507
rect 665 -2473 757 -2467
rect 665 -2507 677 -2473
rect 745 -2507 757 -2473
rect 665 -2513 757 -2507
rect 823 -2473 915 -2467
rect 823 -2507 835 -2473
rect 903 -2507 915 -2473
rect 823 -2513 915 -2507
rect 981 -2473 1073 -2467
rect 981 -2507 993 -2473
rect 1061 -2507 1073 -2473
rect 981 -2513 1073 -2507
rect 1139 -2473 1231 -2467
rect 1139 -2507 1151 -2473
rect 1219 -2507 1231 -2473
rect 1139 -2513 1231 -2507
rect 1297 -2473 1389 -2467
rect 1297 -2507 1309 -2473
rect 1377 -2507 1389 -2473
rect 1297 -2513 1389 -2507
rect 1455 -2473 1547 -2467
rect 1455 -2507 1467 -2473
rect 1535 -2507 1547 -2473
rect 1455 -2513 1547 -2507
rect -1603 -2557 -1557 -2545
rect -1603 -3533 -1597 -2557
rect -1563 -3533 -1557 -2557
rect -1603 -3545 -1557 -3533
rect -1445 -2557 -1399 -2545
rect -1445 -3533 -1439 -2557
rect -1405 -3533 -1399 -2557
rect -1445 -3545 -1399 -3533
rect -1287 -2557 -1241 -2545
rect -1287 -3533 -1281 -2557
rect -1247 -3533 -1241 -2557
rect -1287 -3545 -1241 -3533
rect -1129 -2557 -1083 -2545
rect -1129 -3533 -1123 -2557
rect -1089 -3533 -1083 -2557
rect -1129 -3545 -1083 -3533
rect -971 -2557 -925 -2545
rect -971 -3533 -965 -2557
rect -931 -3533 -925 -2557
rect -971 -3545 -925 -3533
rect -813 -2557 -767 -2545
rect -813 -3533 -807 -2557
rect -773 -3533 -767 -2557
rect -813 -3545 -767 -3533
rect -655 -2557 -609 -2545
rect -655 -3533 -649 -2557
rect -615 -3533 -609 -2557
rect -655 -3545 -609 -3533
rect -497 -2557 -451 -2545
rect -497 -3533 -491 -2557
rect -457 -3533 -451 -2557
rect -497 -3545 -451 -3533
rect -339 -2557 -293 -2545
rect -339 -3533 -333 -2557
rect -299 -3533 -293 -2557
rect -339 -3545 -293 -3533
rect -181 -2557 -135 -2545
rect -181 -3533 -175 -2557
rect -141 -3533 -135 -2557
rect -181 -3545 -135 -3533
rect -23 -2557 23 -2545
rect -23 -3533 -17 -2557
rect 17 -3533 23 -2557
rect -23 -3545 23 -3533
rect 135 -2557 181 -2545
rect 135 -3533 141 -2557
rect 175 -3533 181 -2557
rect 135 -3545 181 -3533
rect 293 -2557 339 -2545
rect 293 -3533 299 -2557
rect 333 -3533 339 -2557
rect 293 -3545 339 -3533
rect 451 -2557 497 -2545
rect 451 -3533 457 -2557
rect 491 -3533 497 -2557
rect 451 -3545 497 -3533
rect 609 -2557 655 -2545
rect 609 -3533 615 -2557
rect 649 -3533 655 -2557
rect 609 -3545 655 -3533
rect 767 -2557 813 -2545
rect 767 -3533 773 -2557
rect 807 -3533 813 -2557
rect 767 -3545 813 -3533
rect 925 -2557 971 -2545
rect 925 -3533 931 -2557
rect 965 -3533 971 -2557
rect 925 -3545 971 -3533
rect 1083 -2557 1129 -2545
rect 1083 -3533 1089 -2557
rect 1123 -3533 1129 -2557
rect 1083 -3545 1129 -3533
rect 1241 -2557 1287 -2545
rect 1241 -3533 1247 -2557
rect 1281 -3533 1287 -2557
rect 1241 -3545 1287 -3533
rect 1399 -2557 1445 -2545
rect 1399 -3533 1405 -2557
rect 1439 -3533 1445 -2557
rect 1399 -3545 1445 -3533
rect 1557 -2557 1603 -2545
rect 1557 -3533 1563 -2557
rect 1597 -3533 1603 -2557
rect 1557 -3545 1603 -3533
rect -1547 -3583 -1455 -3577
rect -1547 -3617 -1535 -3583
rect -1467 -3617 -1455 -3583
rect -1547 -3623 -1455 -3617
rect -1389 -3583 -1297 -3577
rect -1389 -3617 -1377 -3583
rect -1309 -3617 -1297 -3583
rect -1389 -3623 -1297 -3617
rect -1231 -3583 -1139 -3577
rect -1231 -3617 -1219 -3583
rect -1151 -3617 -1139 -3583
rect -1231 -3623 -1139 -3617
rect -1073 -3583 -981 -3577
rect -1073 -3617 -1061 -3583
rect -993 -3617 -981 -3583
rect -1073 -3623 -981 -3617
rect -915 -3583 -823 -3577
rect -915 -3617 -903 -3583
rect -835 -3617 -823 -3583
rect -915 -3623 -823 -3617
rect -757 -3583 -665 -3577
rect -757 -3617 -745 -3583
rect -677 -3617 -665 -3583
rect -757 -3623 -665 -3617
rect -599 -3583 -507 -3577
rect -599 -3617 -587 -3583
rect -519 -3617 -507 -3583
rect -599 -3623 -507 -3617
rect -441 -3583 -349 -3577
rect -441 -3617 -429 -3583
rect -361 -3617 -349 -3583
rect -441 -3623 -349 -3617
rect -283 -3583 -191 -3577
rect -283 -3617 -271 -3583
rect -203 -3617 -191 -3583
rect -283 -3623 -191 -3617
rect -125 -3583 -33 -3577
rect -125 -3617 -113 -3583
rect -45 -3617 -33 -3583
rect -125 -3623 -33 -3617
rect 33 -3583 125 -3577
rect 33 -3617 45 -3583
rect 113 -3617 125 -3583
rect 33 -3623 125 -3617
rect 191 -3583 283 -3577
rect 191 -3617 203 -3583
rect 271 -3617 283 -3583
rect 191 -3623 283 -3617
rect 349 -3583 441 -3577
rect 349 -3617 361 -3583
rect 429 -3617 441 -3583
rect 349 -3623 441 -3617
rect 507 -3583 599 -3577
rect 507 -3617 519 -3583
rect 587 -3617 599 -3583
rect 507 -3623 599 -3617
rect 665 -3583 757 -3577
rect 665 -3617 677 -3583
rect 745 -3617 757 -3583
rect 665 -3623 757 -3617
rect 823 -3583 915 -3577
rect 823 -3617 835 -3583
rect 903 -3617 915 -3583
rect 823 -3623 915 -3617
rect 981 -3583 1073 -3577
rect 981 -3617 993 -3583
rect 1061 -3617 1073 -3583
rect 981 -3623 1073 -3617
rect 1139 -3583 1231 -3577
rect 1139 -3617 1151 -3583
rect 1219 -3617 1231 -3583
rect 1139 -3623 1231 -3617
rect 1297 -3583 1389 -3577
rect 1297 -3617 1309 -3583
rect 1377 -3617 1389 -3583
rect 1297 -3623 1389 -3617
rect 1455 -3583 1547 -3577
rect 1455 -3617 1467 -3583
rect 1535 -3617 1547 -3583
rect 1455 -3623 1547 -3617
rect -1547 -3691 -1455 -3685
rect -1547 -3725 -1535 -3691
rect -1467 -3725 -1455 -3691
rect -1547 -3731 -1455 -3725
rect -1389 -3691 -1297 -3685
rect -1389 -3725 -1377 -3691
rect -1309 -3725 -1297 -3691
rect -1389 -3731 -1297 -3725
rect -1231 -3691 -1139 -3685
rect -1231 -3725 -1219 -3691
rect -1151 -3725 -1139 -3691
rect -1231 -3731 -1139 -3725
rect -1073 -3691 -981 -3685
rect -1073 -3725 -1061 -3691
rect -993 -3725 -981 -3691
rect -1073 -3731 -981 -3725
rect -915 -3691 -823 -3685
rect -915 -3725 -903 -3691
rect -835 -3725 -823 -3691
rect -915 -3731 -823 -3725
rect -757 -3691 -665 -3685
rect -757 -3725 -745 -3691
rect -677 -3725 -665 -3691
rect -757 -3731 -665 -3725
rect -599 -3691 -507 -3685
rect -599 -3725 -587 -3691
rect -519 -3725 -507 -3691
rect -599 -3731 -507 -3725
rect -441 -3691 -349 -3685
rect -441 -3725 -429 -3691
rect -361 -3725 -349 -3691
rect -441 -3731 -349 -3725
rect -283 -3691 -191 -3685
rect -283 -3725 -271 -3691
rect -203 -3725 -191 -3691
rect -283 -3731 -191 -3725
rect -125 -3691 -33 -3685
rect -125 -3725 -113 -3691
rect -45 -3725 -33 -3691
rect -125 -3731 -33 -3725
rect 33 -3691 125 -3685
rect 33 -3725 45 -3691
rect 113 -3725 125 -3691
rect 33 -3731 125 -3725
rect 191 -3691 283 -3685
rect 191 -3725 203 -3691
rect 271 -3725 283 -3691
rect 191 -3731 283 -3725
rect 349 -3691 441 -3685
rect 349 -3725 361 -3691
rect 429 -3725 441 -3691
rect 349 -3731 441 -3725
rect 507 -3691 599 -3685
rect 507 -3725 519 -3691
rect 587 -3725 599 -3691
rect 507 -3731 599 -3725
rect 665 -3691 757 -3685
rect 665 -3725 677 -3691
rect 745 -3725 757 -3691
rect 665 -3731 757 -3725
rect 823 -3691 915 -3685
rect 823 -3725 835 -3691
rect 903 -3725 915 -3691
rect 823 -3731 915 -3725
rect 981 -3691 1073 -3685
rect 981 -3725 993 -3691
rect 1061 -3725 1073 -3691
rect 981 -3731 1073 -3725
rect 1139 -3691 1231 -3685
rect 1139 -3725 1151 -3691
rect 1219 -3725 1231 -3691
rect 1139 -3731 1231 -3725
rect 1297 -3691 1389 -3685
rect 1297 -3725 1309 -3691
rect 1377 -3725 1389 -3691
rect 1297 -3731 1389 -3725
rect 1455 -3691 1547 -3685
rect 1455 -3725 1467 -3691
rect 1535 -3725 1547 -3691
rect 1455 -3731 1547 -3725
rect -1603 -3775 -1557 -3763
rect -1603 -4751 -1597 -3775
rect -1563 -4751 -1557 -3775
rect -1603 -4763 -1557 -4751
rect -1445 -3775 -1399 -3763
rect -1445 -4751 -1439 -3775
rect -1405 -4751 -1399 -3775
rect -1445 -4763 -1399 -4751
rect -1287 -3775 -1241 -3763
rect -1287 -4751 -1281 -3775
rect -1247 -4751 -1241 -3775
rect -1287 -4763 -1241 -4751
rect -1129 -3775 -1083 -3763
rect -1129 -4751 -1123 -3775
rect -1089 -4751 -1083 -3775
rect -1129 -4763 -1083 -4751
rect -971 -3775 -925 -3763
rect -971 -4751 -965 -3775
rect -931 -4751 -925 -3775
rect -971 -4763 -925 -4751
rect -813 -3775 -767 -3763
rect -813 -4751 -807 -3775
rect -773 -4751 -767 -3775
rect -813 -4763 -767 -4751
rect -655 -3775 -609 -3763
rect -655 -4751 -649 -3775
rect -615 -4751 -609 -3775
rect -655 -4763 -609 -4751
rect -497 -3775 -451 -3763
rect -497 -4751 -491 -3775
rect -457 -4751 -451 -3775
rect -497 -4763 -451 -4751
rect -339 -3775 -293 -3763
rect -339 -4751 -333 -3775
rect -299 -4751 -293 -3775
rect -339 -4763 -293 -4751
rect -181 -3775 -135 -3763
rect -181 -4751 -175 -3775
rect -141 -4751 -135 -3775
rect -181 -4763 -135 -4751
rect -23 -3775 23 -3763
rect -23 -4751 -17 -3775
rect 17 -4751 23 -3775
rect -23 -4763 23 -4751
rect 135 -3775 181 -3763
rect 135 -4751 141 -3775
rect 175 -4751 181 -3775
rect 135 -4763 181 -4751
rect 293 -3775 339 -3763
rect 293 -4751 299 -3775
rect 333 -4751 339 -3775
rect 293 -4763 339 -4751
rect 451 -3775 497 -3763
rect 451 -4751 457 -3775
rect 491 -4751 497 -3775
rect 451 -4763 497 -4751
rect 609 -3775 655 -3763
rect 609 -4751 615 -3775
rect 649 -4751 655 -3775
rect 609 -4763 655 -4751
rect 767 -3775 813 -3763
rect 767 -4751 773 -3775
rect 807 -4751 813 -3775
rect 767 -4763 813 -4751
rect 925 -3775 971 -3763
rect 925 -4751 931 -3775
rect 965 -4751 971 -3775
rect 925 -4763 971 -4751
rect 1083 -3775 1129 -3763
rect 1083 -4751 1089 -3775
rect 1123 -4751 1129 -3775
rect 1083 -4763 1129 -4751
rect 1241 -3775 1287 -3763
rect 1241 -4751 1247 -3775
rect 1281 -4751 1287 -3775
rect 1241 -4763 1287 -4751
rect 1399 -3775 1445 -3763
rect 1399 -4751 1405 -3775
rect 1439 -4751 1445 -3775
rect 1399 -4763 1445 -4751
rect 1557 -3775 1603 -3763
rect 1557 -4751 1563 -3775
rect 1597 -4751 1603 -3775
rect 1557 -4763 1603 -4751
rect -1547 -4801 -1455 -4795
rect -1547 -4835 -1535 -4801
rect -1467 -4835 -1455 -4801
rect -1547 -4841 -1455 -4835
rect -1389 -4801 -1297 -4795
rect -1389 -4835 -1377 -4801
rect -1309 -4835 -1297 -4801
rect -1389 -4841 -1297 -4835
rect -1231 -4801 -1139 -4795
rect -1231 -4835 -1219 -4801
rect -1151 -4835 -1139 -4801
rect -1231 -4841 -1139 -4835
rect -1073 -4801 -981 -4795
rect -1073 -4835 -1061 -4801
rect -993 -4835 -981 -4801
rect -1073 -4841 -981 -4835
rect -915 -4801 -823 -4795
rect -915 -4835 -903 -4801
rect -835 -4835 -823 -4801
rect -915 -4841 -823 -4835
rect -757 -4801 -665 -4795
rect -757 -4835 -745 -4801
rect -677 -4835 -665 -4801
rect -757 -4841 -665 -4835
rect -599 -4801 -507 -4795
rect -599 -4835 -587 -4801
rect -519 -4835 -507 -4801
rect -599 -4841 -507 -4835
rect -441 -4801 -349 -4795
rect -441 -4835 -429 -4801
rect -361 -4835 -349 -4801
rect -441 -4841 -349 -4835
rect -283 -4801 -191 -4795
rect -283 -4835 -271 -4801
rect -203 -4835 -191 -4801
rect -283 -4841 -191 -4835
rect -125 -4801 -33 -4795
rect -125 -4835 -113 -4801
rect -45 -4835 -33 -4801
rect -125 -4841 -33 -4835
rect 33 -4801 125 -4795
rect 33 -4835 45 -4801
rect 113 -4835 125 -4801
rect 33 -4841 125 -4835
rect 191 -4801 283 -4795
rect 191 -4835 203 -4801
rect 271 -4835 283 -4801
rect 191 -4841 283 -4835
rect 349 -4801 441 -4795
rect 349 -4835 361 -4801
rect 429 -4835 441 -4801
rect 349 -4841 441 -4835
rect 507 -4801 599 -4795
rect 507 -4835 519 -4801
rect 587 -4835 599 -4801
rect 507 -4841 599 -4835
rect 665 -4801 757 -4795
rect 665 -4835 677 -4801
rect 745 -4835 757 -4801
rect 665 -4841 757 -4835
rect 823 -4801 915 -4795
rect 823 -4835 835 -4801
rect 903 -4835 915 -4801
rect 823 -4841 915 -4835
rect 981 -4801 1073 -4795
rect 981 -4835 993 -4801
rect 1061 -4835 1073 -4801
rect 981 -4841 1073 -4835
rect 1139 -4801 1231 -4795
rect 1139 -4835 1151 -4801
rect 1219 -4835 1231 -4801
rect 1139 -4841 1231 -4835
rect 1297 -4801 1389 -4795
rect 1297 -4835 1309 -4801
rect 1377 -4835 1389 -4801
rect 1297 -4841 1389 -4835
rect 1455 -4801 1547 -4795
rect 1455 -4835 1467 -4801
rect 1535 -4835 1547 -4801
rect 1455 -4841 1547 -4835
rect -1547 -4909 -1455 -4903
rect -1547 -4943 -1535 -4909
rect -1467 -4943 -1455 -4909
rect -1547 -4949 -1455 -4943
rect -1389 -4909 -1297 -4903
rect -1389 -4943 -1377 -4909
rect -1309 -4943 -1297 -4909
rect -1389 -4949 -1297 -4943
rect -1231 -4909 -1139 -4903
rect -1231 -4943 -1219 -4909
rect -1151 -4943 -1139 -4909
rect -1231 -4949 -1139 -4943
rect -1073 -4909 -981 -4903
rect -1073 -4943 -1061 -4909
rect -993 -4943 -981 -4909
rect -1073 -4949 -981 -4943
rect -915 -4909 -823 -4903
rect -915 -4943 -903 -4909
rect -835 -4943 -823 -4909
rect -915 -4949 -823 -4943
rect -757 -4909 -665 -4903
rect -757 -4943 -745 -4909
rect -677 -4943 -665 -4909
rect -757 -4949 -665 -4943
rect -599 -4909 -507 -4903
rect -599 -4943 -587 -4909
rect -519 -4943 -507 -4909
rect -599 -4949 -507 -4943
rect -441 -4909 -349 -4903
rect -441 -4943 -429 -4909
rect -361 -4943 -349 -4909
rect -441 -4949 -349 -4943
rect -283 -4909 -191 -4903
rect -283 -4943 -271 -4909
rect -203 -4943 -191 -4909
rect -283 -4949 -191 -4943
rect -125 -4909 -33 -4903
rect -125 -4943 -113 -4909
rect -45 -4943 -33 -4909
rect -125 -4949 -33 -4943
rect 33 -4909 125 -4903
rect 33 -4943 45 -4909
rect 113 -4943 125 -4909
rect 33 -4949 125 -4943
rect 191 -4909 283 -4903
rect 191 -4943 203 -4909
rect 271 -4943 283 -4909
rect 191 -4949 283 -4943
rect 349 -4909 441 -4903
rect 349 -4943 361 -4909
rect 429 -4943 441 -4909
rect 349 -4949 441 -4943
rect 507 -4909 599 -4903
rect 507 -4943 519 -4909
rect 587 -4943 599 -4909
rect 507 -4949 599 -4943
rect 665 -4909 757 -4903
rect 665 -4943 677 -4909
rect 745 -4943 757 -4909
rect 665 -4949 757 -4943
rect 823 -4909 915 -4903
rect 823 -4943 835 -4909
rect 903 -4943 915 -4909
rect 823 -4949 915 -4943
rect 981 -4909 1073 -4903
rect 981 -4943 993 -4909
rect 1061 -4943 1073 -4909
rect 981 -4949 1073 -4943
rect 1139 -4909 1231 -4903
rect 1139 -4943 1151 -4909
rect 1219 -4943 1231 -4909
rect 1139 -4949 1231 -4943
rect 1297 -4909 1389 -4903
rect 1297 -4943 1309 -4909
rect 1377 -4943 1389 -4909
rect 1297 -4949 1389 -4943
rect 1455 -4909 1547 -4903
rect 1455 -4943 1467 -4909
rect 1535 -4943 1547 -4909
rect 1455 -4949 1547 -4943
rect -1603 -4993 -1557 -4981
rect -1603 -5969 -1597 -4993
rect -1563 -5969 -1557 -4993
rect -1603 -5981 -1557 -5969
rect -1445 -4993 -1399 -4981
rect -1445 -5969 -1439 -4993
rect -1405 -5969 -1399 -4993
rect -1445 -5981 -1399 -5969
rect -1287 -4993 -1241 -4981
rect -1287 -5969 -1281 -4993
rect -1247 -5969 -1241 -4993
rect -1287 -5981 -1241 -5969
rect -1129 -4993 -1083 -4981
rect -1129 -5969 -1123 -4993
rect -1089 -5969 -1083 -4993
rect -1129 -5981 -1083 -5969
rect -971 -4993 -925 -4981
rect -971 -5969 -965 -4993
rect -931 -5969 -925 -4993
rect -971 -5981 -925 -5969
rect -813 -4993 -767 -4981
rect -813 -5969 -807 -4993
rect -773 -5969 -767 -4993
rect -813 -5981 -767 -5969
rect -655 -4993 -609 -4981
rect -655 -5969 -649 -4993
rect -615 -5969 -609 -4993
rect -655 -5981 -609 -5969
rect -497 -4993 -451 -4981
rect -497 -5969 -491 -4993
rect -457 -5969 -451 -4993
rect -497 -5981 -451 -5969
rect -339 -4993 -293 -4981
rect -339 -5969 -333 -4993
rect -299 -5969 -293 -4993
rect -339 -5981 -293 -5969
rect -181 -4993 -135 -4981
rect -181 -5969 -175 -4993
rect -141 -5969 -135 -4993
rect -181 -5981 -135 -5969
rect -23 -4993 23 -4981
rect -23 -5969 -17 -4993
rect 17 -5969 23 -4993
rect -23 -5981 23 -5969
rect 135 -4993 181 -4981
rect 135 -5969 141 -4993
rect 175 -5969 181 -4993
rect 135 -5981 181 -5969
rect 293 -4993 339 -4981
rect 293 -5969 299 -4993
rect 333 -5969 339 -4993
rect 293 -5981 339 -5969
rect 451 -4993 497 -4981
rect 451 -5969 457 -4993
rect 491 -5969 497 -4993
rect 451 -5981 497 -5969
rect 609 -4993 655 -4981
rect 609 -5969 615 -4993
rect 649 -5969 655 -4993
rect 609 -5981 655 -5969
rect 767 -4993 813 -4981
rect 767 -5969 773 -4993
rect 807 -5969 813 -4993
rect 767 -5981 813 -5969
rect 925 -4993 971 -4981
rect 925 -5969 931 -4993
rect 965 -5969 971 -4993
rect 925 -5981 971 -5969
rect 1083 -4993 1129 -4981
rect 1083 -5969 1089 -4993
rect 1123 -5969 1129 -4993
rect 1083 -5981 1129 -5969
rect 1241 -4993 1287 -4981
rect 1241 -5969 1247 -4993
rect 1281 -5969 1287 -4993
rect 1241 -5981 1287 -5969
rect 1399 -4993 1445 -4981
rect 1399 -5969 1405 -4993
rect 1439 -5969 1445 -4993
rect 1399 -5981 1445 -5969
rect 1557 -4993 1603 -4981
rect 1557 -5969 1563 -4993
rect 1597 -5969 1603 -4993
rect 1557 -5981 1603 -5969
rect -1547 -6019 -1455 -6013
rect -1547 -6053 -1535 -6019
rect -1467 -6053 -1455 -6019
rect -1547 -6059 -1455 -6053
rect -1389 -6019 -1297 -6013
rect -1389 -6053 -1377 -6019
rect -1309 -6053 -1297 -6019
rect -1389 -6059 -1297 -6053
rect -1231 -6019 -1139 -6013
rect -1231 -6053 -1219 -6019
rect -1151 -6053 -1139 -6019
rect -1231 -6059 -1139 -6053
rect -1073 -6019 -981 -6013
rect -1073 -6053 -1061 -6019
rect -993 -6053 -981 -6019
rect -1073 -6059 -981 -6053
rect -915 -6019 -823 -6013
rect -915 -6053 -903 -6019
rect -835 -6053 -823 -6019
rect -915 -6059 -823 -6053
rect -757 -6019 -665 -6013
rect -757 -6053 -745 -6019
rect -677 -6053 -665 -6019
rect -757 -6059 -665 -6053
rect -599 -6019 -507 -6013
rect -599 -6053 -587 -6019
rect -519 -6053 -507 -6019
rect -599 -6059 -507 -6053
rect -441 -6019 -349 -6013
rect -441 -6053 -429 -6019
rect -361 -6053 -349 -6019
rect -441 -6059 -349 -6053
rect -283 -6019 -191 -6013
rect -283 -6053 -271 -6019
rect -203 -6053 -191 -6019
rect -283 -6059 -191 -6053
rect -125 -6019 -33 -6013
rect -125 -6053 -113 -6019
rect -45 -6053 -33 -6019
rect -125 -6059 -33 -6053
rect 33 -6019 125 -6013
rect 33 -6053 45 -6019
rect 113 -6053 125 -6019
rect 33 -6059 125 -6053
rect 191 -6019 283 -6013
rect 191 -6053 203 -6019
rect 271 -6053 283 -6019
rect 191 -6059 283 -6053
rect 349 -6019 441 -6013
rect 349 -6053 361 -6019
rect 429 -6053 441 -6019
rect 349 -6059 441 -6053
rect 507 -6019 599 -6013
rect 507 -6053 519 -6019
rect 587 -6053 599 -6019
rect 507 -6059 599 -6053
rect 665 -6019 757 -6013
rect 665 -6053 677 -6019
rect 745 -6053 757 -6019
rect 665 -6059 757 -6053
rect 823 -6019 915 -6013
rect 823 -6053 835 -6019
rect 903 -6053 915 -6019
rect 823 -6059 915 -6053
rect 981 -6019 1073 -6013
rect 981 -6053 993 -6019
rect 1061 -6053 1073 -6019
rect 981 -6059 1073 -6053
rect 1139 -6019 1231 -6013
rect 1139 -6053 1151 -6019
rect 1219 -6053 1231 -6019
rect 1139 -6059 1231 -6053
rect 1297 -6019 1389 -6013
rect 1297 -6053 1309 -6019
rect 1377 -6053 1389 -6019
rect 1297 -6059 1389 -6053
rect 1455 -6019 1547 -6013
rect 1455 -6053 1467 -6019
rect 1535 -6053 1547 -6019
rect 1455 -6059 1547 -6053
<< properties >>
string FIXED_BBOX -1714 -6174 1714 6174
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string MASKHINTS_HVI -1790 -6240 1790 6240
string parameters w 5.0 l 0.5 m 10 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
