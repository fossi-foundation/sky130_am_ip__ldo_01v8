magic
tech sky130A
magscale 1 2
timestamp 1717294357
<< metal3 >>
rect -686 512 686 540
rect -686 -512 602 512
rect 666 -512 686 512
rect -686 -540 686 -512
<< via3 >>
rect 602 -512 666 512
<< mimcap >>
rect -646 460 354 500
rect -646 -460 -606 460
rect 314 -460 354 460
rect -646 -500 354 -460
<< mimcapcontact >>
rect -606 -460 314 460
<< metal4 >>
rect 586 512 682 528
rect -607 460 315 461
rect -607 -460 -606 460
rect 314 -460 315 460
rect -607 -461 315 -460
rect 586 -512 602 512
rect 666 -512 682 512
rect 586 -528 682 -512
<< properties >>
string FIXED_BBOX -686 -540 394 540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
