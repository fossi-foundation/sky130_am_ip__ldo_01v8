magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< pwell >>
rect -278 -1403 278 1403
<< mvnmos >>
rect -50 945 50 1145
rect -50 527 50 727
rect -50 109 50 309
rect -50 -309 50 -109
rect -50 -727 50 -527
rect -50 -1145 50 -945
<< mvndiff >>
rect -108 1133 -50 1145
rect -108 957 -96 1133
rect -62 957 -50 1133
rect -108 945 -50 957
rect 50 1133 108 1145
rect 50 957 62 1133
rect 96 957 108 1133
rect 50 945 108 957
rect -108 715 -50 727
rect -108 539 -96 715
rect -62 539 -50 715
rect -108 527 -50 539
rect 50 715 108 727
rect 50 539 62 715
rect 96 539 108 715
rect 50 527 108 539
rect -108 297 -50 309
rect -108 121 -96 297
rect -62 121 -50 297
rect -108 109 -50 121
rect 50 297 108 309
rect 50 121 62 297
rect 96 121 108 297
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -297 -96 -121
rect -62 -297 -50 -121
rect -108 -309 -50 -297
rect 50 -121 108 -109
rect 50 -297 62 -121
rect 96 -297 108 -121
rect 50 -309 108 -297
rect -108 -539 -50 -527
rect -108 -715 -96 -539
rect -62 -715 -50 -539
rect -108 -727 -50 -715
rect 50 -539 108 -527
rect 50 -715 62 -539
rect 96 -715 108 -539
rect 50 -727 108 -715
rect -108 -957 -50 -945
rect -108 -1133 -96 -957
rect -62 -1133 -50 -957
rect -108 -1145 -50 -1133
rect 50 -957 108 -945
rect 50 -1133 62 -957
rect 96 -1133 108 -957
rect 50 -1145 108 -1133
<< mvndiffc >>
rect -96 957 -62 1133
rect 62 957 96 1133
rect -96 539 -62 715
rect 62 539 96 715
rect -96 121 -62 297
rect 62 121 96 297
rect -96 -297 -62 -121
rect 62 -297 96 -121
rect -96 -715 -62 -539
rect 62 -715 96 -539
rect -96 -1133 -62 -957
rect 62 -1133 96 -957
<< mvpsubdiff >>
rect -242 1355 242 1367
rect -242 1321 -134 1355
rect 134 1321 242 1355
rect -242 1309 242 1321
rect -242 1259 -184 1309
rect -242 -1259 -230 1259
rect -196 -1259 -184 1259
rect 184 1259 242 1309
rect -242 -1309 -184 -1259
rect 184 -1259 196 1259
rect 230 -1259 242 1259
rect 184 -1309 242 -1259
rect -242 -1321 242 -1309
rect -242 -1355 -134 -1321
rect 134 -1355 242 -1321
rect -242 -1367 242 -1355
<< mvpsubdiffcont >>
rect -134 1321 134 1355
rect -230 -1259 -196 1259
rect 196 -1259 230 1259
rect -134 -1355 134 -1321
<< poly >>
rect -50 1217 50 1233
rect -50 1183 -34 1217
rect 34 1183 50 1217
rect -50 1145 50 1183
rect -50 907 50 945
rect -50 873 -34 907
rect 34 873 50 907
rect -50 857 50 873
rect -50 799 50 815
rect -50 765 -34 799
rect 34 765 50 799
rect -50 727 50 765
rect -50 489 50 527
rect -50 455 -34 489
rect 34 455 50 489
rect -50 439 50 455
rect -50 381 50 397
rect -50 347 -34 381
rect 34 347 50 381
rect -50 309 50 347
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -347 50 -309
rect -50 -381 -34 -347
rect 34 -381 50 -347
rect -50 -397 50 -381
rect -50 -455 50 -439
rect -50 -489 -34 -455
rect 34 -489 50 -455
rect -50 -527 50 -489
rect -50 -765 50 -727
rect -50 -799 -34 -765
rect 34 -799 50 -765
rect -50 -815 50 -799
rect -50 -873 50 -857
rect -50 -907 -34 -873
rect 34 -907 50 -873
rect -50 -945 50 -907
rect -50 -1183 50 -1145
rect -50 -1217 -34 -1183
rect 34 -1217 50 -1183
rect -50 -1233 50 -1217
<< polycont >>
rect -34 1183 34 1217
rect -34 873 34 907
rect -34 765 34 799
rect -34 455 34 489
rect -34 347 34 381
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -381 34 -347
rect -34 -489 34 -455
rect -34 -799 34 -765
rect -34 -907 34 -873
rect -34 -1217 34 -1183
<< locali >>
rect -230 1321 -134 1355
rect 134 1321 230 1355
rect -230 1259 -196 1321
rect 196 1259 230 1321
rect -50 1183 -34 1217
rect 34 1183 50 1217
rect -96 1133 -62 1149
rect -96 941 -62 957
rect 62 1133 96 1149
rect 62 941 96 957
rect -50 873 -34 907
rect 34 873 50 907
rect -50 765 -34 799
rect 34 765 50 799
rect -96 715 -62 731
rect -96 523 -62 539
rect 62 715 96 731
rect 62 523 96 539
rect -50 455 -34 489
rect 34 455 50 489
rect -50 347 -34 381
rect 34 347 50 381
rect -96 297 -62 313
rect -96 105 -62 121
rect 62 297 96 313
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -313 -62 -297
rect 62 -121 96 -105
rect 62 -313 96 -297
rect -50 -381 -34 -347
rect 34 -381 50 -347
rect -50 -489 -34 -455
rect 34 -489 50 -455
rect -96 -539 -62 -523
rect -96 -731 -62 -715
rect 62 -539 96 -523
rect 62 -731 96 -715
rect -50 -799 -34 -765
rect 34 -799 50 -765
rect -50 -907 -34 -873
rect 34 -907 50 -873
rect -96 -957 -62 -941
rect -96 -1149 -62 -1133
rect 62 -957 96 -941
rect 62 -1149 96 -1133
rect -50 -1217 -34 -1183
rect 34 -1217 50 -1183
rect -230 -1321 -196 -1259
rect 196 -1321 230 -1259
rect -230 -1355 -134 -1321
rect 134 -1355 230 -1321
<< viali >>
rect -34 1183 34 1217
rect -96 957 -62 1133
rect 62 957 96 1133
rect -34 873 34 907
rect -34 765 34 799
rect -96 539 -62 715
rect 62 539 96 715
rect -34 455 34 489
rect -34 347 34 381
rect -96 121 -62 297
rect 62 121 96 297
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -297 -62 -121
rect 62 -297 96 -121
rect -34 -381 34 -347
rect -34 -489 34 -455
rect -96 -715 -62 -539
rect 62 -715 96 -539
rect -34 -799 34 -765
rect -34 -907 34 -873
rect -96 -1133 -62 -957
rect 62 -1133 96 -957
rect -34 -1217 34 -1183
<< metal1 >>
rect -46 1217 46 1223
rect -46 1183 -34 1217
rect 34 1183 46 1217
rect -46 1177 46 1183
rect -102 1133 -56 1145
rect -102 957 -96 1133
rect -62 957 -56 1133
rect -102 945 -56 957
rect 56 1133 102 1145
rect 56 957 62 1133
rect 96 957 102 1133
rect 56 945 102 957
rect -46 907 46 913
rect -46 873 -34 907
rect 34 873 46 907
rect -46 867 46 873
rect -46 799 46 805
rect -46 765 -34 799
rect 34 765 46 799
rect -46 759 46 765
rect -102 715 -56 727
rect -102 539 -96 715
rect -62 539 -56 715
rect -102 527 -56 539
rect 56 715 102 727
rect 56 539 62 715
rect 96 539 102 715
rect 56 527 102 539
rect -46 489 46 495
rect -46 455 -34 489
rect 34 455 46 489
rect -46 449 46 455
rect -46 381 46 387
rect -46 347 -34 381
rect 34 347 46 381
rect -46 341 46 347
rect -102 297 -56 309
rect -102 121 -96 297
rect -62 121 -56 297
rect -102 109 -56 121
rect 56 297 102 309
rect 56 121 62 297
rect 96 121 102 297
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -297 -96 -121
rect -62 -297 -56 -121
rect -102 -309 -56 -297
rect 56 -121 102 -109
rect 56 -297 62 -121
rect 96 -297 102 -121
rect 56 -309 102 -297
rect -46 -347 46 -341
rect -46 -381 -34 -347
rect 34 -381 46 -347
rect -46 -387 46 -381
rect -46 -455 46 -449
rect -46 -489 -34 -455
rect 34 -489 46 -455
rect -46 -495 46 -489
rect -102 -539 -56 -527
rect -102 -715 -96 -539
rect -62 -715 -56 -539
rect -102 -727 -56 -715
rect 56 -539 102 -527
rect 56 -715 62 -539
rect 96 -715 102 -539
rect 56 -727 102 -715
rect -46 -765 46 -759
rect -46 -799 -34 -765
rect 34 -799 46 -765
rect -46 -805 46 -799
rect -46 -873 46 -867
rect -46 -907 -34 -873
rect 34 -907 46 -873
rect -46 -913 46 -907
rect -102 -957 -56 -945
rect -102 -1133 -96 -957
rect -62 -1133 -56 -957
rect -102 -1145 -56 -1133
rect 56 -957 102 -945
rect 56 -1133 62 -957
rect 96 -1133 102 -957
rect 56 -1145 102 -1133
rect -46 -1183 46 -1177
rect -46 -1217 -34 -1183
rect 34 -1217 46 -1183
rect -46 -1223 46 -1217
<< properties >>
string FIXED_BBOX -213 -1338 213 1338
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
