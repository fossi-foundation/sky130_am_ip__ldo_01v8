magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -1258 -2359 1258 2359
<< mvpmos >>
rect -1000 1862 1000 2062
rect -1000 1426 1000 1626
rect -1000 990 1000 1190
rect -1000 554 1000 754
rect -1000 118 1000 318
rect -1000 -318 1000 -118
rect -1000 -754 1000 -554
rect -1000 -1190 1000 -990
rect -1000 -1626 1000 -1426
rect -1000 -2062 1000 -1862
<< mvpdiff >>
rect -1058 2050 -1000 2062
rect -1058 1874 -1046 2050
rect -1012 1874 -1000 2050
rect -1058 1862 -1000 1874
rect 1000 2050 1058 2062
rect 1000 1874 1012 2050
rect 1046 1874 1058 2050
rect 1000 1862 1058 1874
rect -1058 1614 -1000 1626
rect -1058 1438 -1046 1614
rect -1012 1438 -1000 1614
rect -1058 1426 -1000 1438
rect 1000 1614 1058 1626
rect 1000 1438 1012 1614
rect 1046 1438 1058 1614
rect 1000 1426 1058 1438
rect -1058 1178 -1000 1190
rect -1058 1002 -1046 1178
rect -1012 1002 -1000 1178
rect -1058 990 -1000 1002
rect 1000 1178 1058 1190
rect 1000 1002 1012 1178
rect 1046 1002 1058 1178
rect 1000 990 1058 1002
rect -1058 742 -1000 754
rect -1058 566 -1046 742
rect -1012 566 -1000 742
rect -1058 554 -1000 566
rect 1000 742 1058 754
rect 1000 566 1012 742
rect 1046 566 1058 742
rect 1000 554 1058 566
rect -1058 306 -1000 318
rect -1058 130 -1046 306
rect -1012 130 -1000 306
rect -1058 118 -1000 130
rect 1000 306 1058 318
rect 1000 130 1012 306
rect 1046 130 1058 306
rect 1000 118 1058 130
rect -1058 -130 -1000 -118
rect -1058 -306 -1046 -130
rect -1012 -306 -1000 -130
rect -1058 -318 -1000 -306
rect 1000 -130 1058 -118
rect 1000 -306 1012 -130
rect 1046 -306 1058 -130
rect 1000 -318 1058 -306
rect -1058 -566 -1000 -554
rect -1058 -742 -1046 -566
rect -1012 -742 -1000 -566
rect -1058 -754 -1000 -742
rect 1000 -566 1058 -554
rect 1000 -742 1012 -566
rect 1046 -742 1058 -566
rect 1000 -754 1058 -742
rect -1058 -1002 -1000 -990
rect -1058 -1178 -1046 -1002
rect -1012 -1178 -1000 -1002
rect -1058 -1190 -1000 -1178
rect 1000 -1002 1058 -990
rect 1000 -1178 1012 -1002
rect 1046 -1178 1058 -1002
rect 1000 -1190 1058 -1178
rect -1058 -1438 -1000 -1426
rect -1058 -1614 -1046 -1438
rect -1012 -1614 -1000 -1438
rect -1058 -1626 -1000 -1614
rect 1000 -1438 1058 -1426
rect 1000 -1614 1012 -1438
rect 1046 -1614 1058 -1438
rect 1000 -1626 1058 -1614
rect -1058 -1874 -1000 -1862
rect -1058 -2050 -1046 -1874
rect -1012 -2050 -1000 -1874
rect -1058 -2062 -1000 -2050
rect 1000 -1874 1058 -1862
rect 1000 -2050 1012 -1874
rect 1046 -2050 1058 -1874
rect 1000 -2062 1058 -2050
<< mvpdiffc >>
rect -1046 1874 -1012 2050
rect 1012 1874 1046 2050
rect -1046 1438 -1012 1614
rect 1012 1438 1046 1614
rect -1046 1002 -1012 1178
rect 1012 1002 1046 1178
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
rect -1046 -1178 -1012 -1002
rect 1012 -1178 1046 -1002
rect -1046 -1614 -1012 -1438
rect 1012 -1614 1046 -1438
rect -1046 -2050 -1012 -1874
rect 1012 -2050 1046 -1874
<< mvnsubdiff >>
rect -1192 2281 1192 2293
rect -1192 2247 -1084 2281
rect 1084 2247 1192 2281
rect -1192 2235 1192 2247
rect -1192 2185 -1134 2235
rect -1192 -2185 -1180 2185
rect -1146 -2185 -1134 2185
rect 1134 2185 1192 2235
rect -1192 -2235 -1134 -2185
rect 1134 -2185 1146 2185
rect 1180 -2185 1192 2185
rect 1134 -2235 1192 -2185
rect -1192 -2247 1192 -2235
rect -1192 -2281 -1084 -2247
rect 1084 -2281 1192 -2247
rect -1192 -2293 1192 -2281
<< mvnsubdiffcont >>
rect -1084 2247 1084 2281
rect -1180 -2185 -1146 2185
rect 1146 -2185 1180 2185
rect -1084 -2281 1084 -2247
<< poly >>
rect -1000 2143 1000 2159
rect -1000 2109 -984 2143
rect 984 2109 1000 2143
rect -1000 2062 1000 2109
rect -1000 1815 1000 1862
rect -1000 1781 -984 1815
rect 984 1781 1000 1815
rect -1000 1765 1000 1781
rect -1000 1707 1000 1723
rect -1000 1673 -984 1707
rect 984 1673 1000 1707
rect -1000 1626 1000 1673
rect -1000 1379 1000 1426
rect -1000 1345 -984 1379
rect 984 1345 1000 1379
rect -1000 1329 1000 1345
rect -1000 1271 1000 1287
rect -1000 1237 -984 1271
rect 984 1237 1000 1271
rect -1000 1190 1000 1237
rect -1000 943 1000 990
rect -1000 909 -984 943
rect 984 909 1000 943
rect -1000 893 1000 909
rect -1000 835 1000 851
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1000 754 1000 801
rect -1000 507 1000 554
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 457 1000 473
rect -1000 399 1000 415
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1000 318 1000 365
rect -1000 71 1000 118
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -118 1000 -71
rect -1000 -365 1000 -318
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -415 1000 -399
rect -1000 -473 1000 -457
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1000 -554 1000 -507
rect -1000 -801 1000 -754
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect -1000 -851 1000 -835
rect -1000 -909 1000 -893
rect -1000 -943 -984 -909
rect 984 -943 1000 -909
rect -1000 -990 1000 -943
rect -1000 -1237 1000 -1190
rect -1000 -1271 -984 -1237
rect 984 -1271 1000 -1237
rect -1000 -1287 1000 -1271
rect -1000 -1345 1000 -1329
rect -1000 -1379 -984 -1345
rect 984 -1379 1000 -1345
rect -1000 -1426 1000 -1379
rect -1000 -1673 1000 -1626
rect -1000 -1707 -984 -1673
rect 984 -1707 1000 -1673
rect -1000 -1723 1000 -1707
rect -1000 -1781 1000 -1765
rect -1000 -1815 -984 -1781
rect 984 -1815 1000 -1781
rect -1000 -1862 1000 -1815
rect -1000 -2109 1000 -2062
rect -1000 -2143 -984 -2109
rect 984 -2143 1000 -2109
rect -1000 -2159 1000 -2143
<< polycont >>
rect -984 2109 984 2143
rect -984 1781 984 1815
rect -984 1673 984 1707
rect -984 1345 984 1379
rect -984 1237 984 1271
rect -984 909 984 943
rect -984 801 984 835
rect -984 473 984 507
rect -984 365 984 399
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -399 984 -365
rect -984 -507 984 -473
rect -984 -835 984 -801
rect -984 -943 984 -909
rect -984 -1271 984 -1237
rect -984 -1379 984 -1345
rect -984 -1707 984 -1673
rect -984 -1815 984 -1781
rect -984 -2143 984 -2109
<< locali >>
rect -1180 2247 -1084 2281
rect 1084 2247 1180 2281
rect -1180 2185 -1146 2247
rect 1146 2185 1180 2247
rect -1000 2109 -984 2143
rect 984 2109 1000 2143
rect -1046 2050 -1012 2066
rect -1046 1858 -1012 1874
rect 1012 2050 1046 2066
rect 1012 1858 1046 1874
rect -1000 1781 -984 1815
rect 984 1781 1000 1815
rect -1000 1673 -984 1707
rect 984 1673 1000 1707
rect -1046 1614 -1012 1630
rect -1046 1422 -1012 1438
rect 1012 1614 1046 1630
rect 1012 1422 1046 1438
rect -1000 1345 -984 1379
rect 984 1345 1000 1379
rect -1000 1237 -984 1271
rect 984 1237 1000 1271
rect -1046 1178 -1012 1194
rect -1046 986 -1012 1002
rect 1012 1178 1046 1194
rect 1012 986 1046 1002
rect -1000 909 -984 943
rect 984 909 1000 943
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1046 742 -1012 758
rect -1046 550 -1012 566
rect 1012 742 1046 758
rect 1012 550 1046 566
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1046 306 -1012 322
rect -1046 114 -1012 130
rect 1012 306 1046 322
rect 1012 114 1046 130
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -130 -1012 -114
rect -1046 -322 -1012 -306
rect 1012 -130 1046 -114
rect 1012 -322 1046 -306
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1046 -566 -1012 -550
rect -1046 -758 -1012 -742
rect 1012 -566 1046 -550
rect 1012 -758 1046 -742
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect -1000 -943 -984 -909
rect 984 -943 1000 -909
rect -1046 -1002 -1012 -986
rect -1046 -1194 -1012 -1178
rect 1012 -1002 1046 -986
rect 1012 -1194 1046 -1178
rect -1000 -1271 -984 -1237
rect 984 -1271 1000 -1237
rect -1000 -1379 -984 -1345
rect 984 -1379 1000 -1345
rect -1046 -1438 -1012 -1422
rect -1046 -1630 -1012 -1614
rect 1012 -1438 1046 -1422
rect 1012 -1630 1046 -1614
rect -1000 -1707 -984 -1673
rect 984 -1707 1000 -1673
rect -1000 -1815 -984 -1781
rect 984 -1815 1000 -1781
rect -1046 -1874 -1012 -1858
rect -1046 -2066 -1012 -2050
rect 1012 -1874 1046 -1858
rect 1012 -2066 1046 -2050
rect -1000 -2143 -984 -2109
rect 984 -2143 1000 -2109
rect -1180 -2247 -1146 -2185
rect 1146 -2247 1180 -2185
rect -1180 -2281 -1084 -2247
rect 1084 -2281 1180 -2247
<< viali >>
rect -984 2109 984 2143
rect -1046 1874 -1012 2050
rect 1012 1874 1046 2050
rect -984 1781 984 1815
rect -984 1673 984 1707
rect -1046 1438 -1012 1614
rect 1012 1438 1046 1614
rect -984 1345 984 1379
rect -984 1237 984 1271
rect -1046 1002 -1012 1178
rect 1012 1002 1046 1178
rect -984 909 984 943
rect -984 801 984 835
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -984 473 984 507
rect -984 365 984 399
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -984 -399 984 -365
rect -984 -507 984 -473
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
rect -984 -835 984 -801
rect -984 -943 984 -909
rect -1046 -1178 -1012 -1002
rect 1012 -1178 1046 -1002
rect -984 -1271 984 -1237
rect -984 -1379 984 -1345
rect -1046 -1614 -1012 -1438
rect 1012 -1614 1046 -1438
rect -984 -1707 984 -1673
rect -984 -1815 984 -1781
rect -1046 -2050 -1012 -1874
rect 1012 -2050 1046 -1874
rect -984 -2143 984 -2109
<< metal1 >>
rect -996 2143 996 2149
rect -996 2109 -984 2143
rect 984 2109 996 2143
rect -996 2103 996 2109
rect -1052 2050 -1006 2062
rect -1052 1874 -1046 2050
rect -1012 1874 -1006 2050
rect -1052 1862 -1006 1874
rect 1006 2050 1052 2062
rect 1006 1874 1012 2050
rect 1046 1874 1052 2050
rect 1006 1862 1052 1874
rect -996 1815 996 1821
rect -996 1781 -984 1815
rect 984 1781 996 1815
rect -996 1775 996 1781
rect -996 1707 996 1713
rect -996 1673 -984 1707
rect 984 1673 996 1707
rect -996 1667 996 1673
rect -1052 1614 -1006 1626
rect -1052 1438 -1046 1614
rect -1012 1438 -1006 1614
rect -1052 1426 -1006 1438
rect 1006 1614 1052 1626
rect 1006 1438 1012 1614
rect 1046 1438 1052 1614
rect 1006 1426 1052 1438
rect -996 1379 996 1385
rect -996 1345 -984 1379
rect 984 1345 996 1379
rect -996 1339 996 1345
rect -996 1271 996 1277
rect -996 1237 -984 1271
rect 984 1237 996 1271
rect -996 1231 996 1237
rect -1052 1178 -1006 1190
rect -1052 1002 -1046 1178
rect -1012 1002 -1006 1178
rect -1052 990 -1006 1002
rect 1006 1178 1052 1190
rect 1006 1002 1012 1178
rect 1046 1002 1052 1178
rect 1006 990 1052 1002
rect -996 943 996 949
rect -996 909 -984 943
rect 984 909 996 943
rect -996 903 996 909
rect -996 835 996 841
rect -996 801 -984 835
rect 984 801 996 835
rect -996 795 996 801
rect -1052 742 -1006 754
rect -1052 566 -1046 742
rect -1012 566 -1006 742
rect -1052 554 -1006 566
rect 1006 742 1052 754
rect 1006 566 1012 742
rect 1046 566 1052 742
rect 1006 554 1052 566
rect -996 507 996 513
rect -996 473 -984 507
rect 984 473 996 507
rect -996 467 996 473
rect -996 399 996 405
rect -996 365 -984 399
rect 984 365 996 399
rect -996 359 996 365
rect -1052 306 -1006 318
rect -1052 130 -1046 306
rect -1012 130 -1006 306
rect -1052 118 -1006 130
rect 1006 306 1052 318
rect 1006 130 1012 306
rect 1046 130 1052 306
rect 1006 118 1052 130
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -130 -1006 -118
rect -1052 -306 -1046 -130
rect -1012 -306 -1006 -130
rect -1052 -318 -1006 -306
rect 1006 -130 1052 -118
rect 1006 -306 1012 -130
rect 1046 -306 1052 -130
rect 1006 -318 1052 -306
rect -996 -365 996 -359
rect -996 -399 -984 -365
rect 984 -399 996 -365
rect -996 -405 996 -399
rect -996 -473 996 -467
rect -996 -507 -984 -473
rect 984 -507 996 -473
rect -996 -513 996 -507
rect -1052 -566 -1006 -554
rect -1052 -742 -1046 -566
rect -1012 -742 -1006 -566
rect -1052 -754 -1006 -742
rect 1006 -566 1052 -554
rect 1006 -742 1012 -566
rect 1046 -742 1052 -566
rect 1006 -754 1052 -742
rect -996 -801 996 -795
rect -996 -835 -984 -801
rect 984 -835 996 -801
rect -996 -841 996 -835
rect -996 -909 996 -903
rect -996 -943 -984 -909
rect 984 -943 996 -909
rect -996 -949 996 -943
rect -1052 -1002 -1006 -990
rect -1052 -1178 -1046 -1002
rect -1012 -1178 -1006 -1002
rect -1052 -1190 -1006 -1178
rect 1006 -1002 1052 -990
rect 1006 -1178 1012 -1002
rect 1046 -1178 1052 -1002
rect 1006 -1190 1052 -1178
rect -996 -1237 996 -1231
rect -996 -1271 -984 -1237
rect 984 -1271 996 -1237
rect -996 -1277 996 -1271
rect -996 -1345 996 -1339
rect -996 -1379 -984 -1345
rect 984 -1379 996 -1345
rect -996 -1385 996 -1379
rect -1052 -1438 -1006 -1426
rect -1052 -1614 -1046 -1438
rect -1012 -1614 -1006 -1438
rect -1052 -1626 -1006 -1614
rect 1006 -1438 1052 -1426
rect 1006 -1614 1012 -1438
rect 1046 -1614 1052 -1438
rect 1006 -1626 1052 -1614
rect -996 -1673 996 -1667
rect -996 -1707 -984 -1673
rect 984 -1707 996 -1673
rect -996 -1713 996 -1707
rect -996 -1781 996 -1775
rect -996 -1815 -984 -1781
rect 984 -1815 996 -1781
rect -996 -1821 996 -1815
rect -1052 -1874 -1006 -1862
rect -1052 -2050 -1046 -1874
rect -1012 -2050 -1006 -1874
rect -1052 -2062 -1006 -2050
rect 1006 -1874 1052 -1862
rect 1006 -2050 1012 -1874
rect 1046 -2050 1052 -1874
rect 1006 -2062 1052 -2050
rect -996 -2109 996 -2103
rect -996 -2143 -984 -2109
rect 984 -2143 996 -2109
rect -996 -2149 996 -2143
<< properties >>
string FIXED_BBOX -1163 -2264 1163 2264
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
