magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -308 -647 308 647
<< mvpmos >>
rect -50 -350 50 350
<< mvpdiff >>
rect -108 338 -50 350
rect -108 -338 -96 338
rect -62 -338 -50 338
rect -108 -350 -50 -338
rect 50 338 108 350
rect 50 -338 62 338
rect 96 -338 108 338
rect 50 -350 108 -338
<< mvpdiffc >>
rect -96 -338 -62 338
rect 62 -338 96 338
<< mvnsubdiff >>
rect -242 569 242 581
rect -242 535 -134 569
rect 134 535 242 569
rect -242 523 242 535
rect -242 473 -184 523
rect -242 -473 -230 473
rect -196 -473 -184 473
rect 184 473 242 523
rect -242 -523 -184 -473
rect 184 -473 196 473
rect 230 -473 242 473
rect 184 -523 242 -473
rect -242 -535 242 -523
rect -242 -569 -134 -535
rect 134 -569 242 -535
rect -242 -581 242 -569
<< mvnsubdiffcont >>
rect -134 535 134 569
rect -230 -473 -196 473
rect 196 -473 230 473
rect -134 -569 134 -535
<< poly >>
rect -50 431 50 447
rect -50 397 -34 431
rect 34 397 50 431
rect -50 350 50 397
rect -50 -397 50 -350
rect -50 -431 -34 -397
rect 34 -431 50 -397
rect -50 -447 50 -431
<< polycont >>
rect -34 397 34 431
rect -34 -431 34 -397
<< locali >>
rect -230 535 -134 569
rect 134 535 230 569
rect -230 473 -196 535
rect 196 473 230 535
rect -50 397 -34 431
rect 34 397 50 431
rect -96 338 -62 354
rect -96 -354 -62 -338
rect 62 338 96 354
rect 62 -354 96 -338
rect -50 -431 -34 -397
rect 34 -431 50 -397
rect -230 -535 -196 -473
rect 196 -535 230 -473
rect -230 -569 -134 -535
rect 134 -569 230 -535
<< viali >>
rect -34 397 34 431
rect -96 -338 -62 338
rect 62 -338 96 338
rect -34 -431 34 -397
<< metal1 >>
rect -46 431 46 437
rect -46 397 -34 431
rect 34 397 46 431
rect -46 391 46 397
rect -102 338 -56 350
rect -102 -338 -96 338
rect -62 -338 -56 338
rect -102 -350 -56 -338
rect 56 338 102 350
rect 56 -338 62 338
rect 96 -338 102 338
rect 56 -350 102 -338
rect -46 -397 46 -391
rect -46 -431 -34 -397
rect 34 -431 46 -397
rect -46 -437 46 -431
<< properties >>
string FIXED_BBOX -213 -552 213 552
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
