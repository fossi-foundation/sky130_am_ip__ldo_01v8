magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< pwell >>
rect -1228 -567 1228 567
<< mvnmos >>
rect -1000 109 1000 309
rect -1000 -309 1000 -109
<< mvndiff >>
rect -1058 297 -1000 309
rect -1058 121 -1046 297
rect -1012 121 -1000 297
rect -1058 109 -1000 121
rect 1000 297 1058 309
rect 1000 121 1012 297
rect 1046 121 1058 297
rect 1000 109 1058 121
rect -1058 -121 -1000 -109
rect -1058 -297 -1046 -121
rect -1012 -297 -1000 -121
rect -1058 -309 -1000 -297
rect 1000 -121 1058 -109
rect 1000 -297 1012 -121
rect 1046 -297 1058 -121
rect 1000 -309 1058 -297
<< mvndiffc >>
rect -1046 121 -1012 297
rect 1012 121 1046 297
rect -1046 -297 -1012 -121
rect 1012 -297 1046 -121
<< mvpsubdiff >>
rect -1192 519 1192 531
rect -1192 485 -1084 519
rect 1084 485 1192 519
rect -1192 473 1192 485
rect -1192 423 -1134 473
rect -1192 -423 -1180 423
rect -1146 -423 -1134 423
rect 1134 423 1192 473
rect -1192 -473 -1134 -423
rect 1134 -423 1146 423
rect 1180 -423 1192 423
rect 1134 -473 1192 -423
rect -1192 -485 1192 -473
rect -1192 -519 -1084 -485
rect 1084 -519 1192 -485
rect -1192 -531 1192 -519
<< mvpsubdiffcont >>
rect -1084 485 1084 519
rect -1180 -423 -1146 423
rect 1146 -423 1180 423
rect -1084 -519 1084 -485
<< poly >>
rect -1000 381 1000 397
rect -1000 347 -984 381
rect 984 347 1000 381
rect -1000 309 1000 347
rect -1000 71 1000 109
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -109 1000 -71
rect -1000 -347 1000 -309
rect -1000 -381 -984 -347
rect 984 -381 1000 -347
rect -1000 -397 1000 -381
<< polycont >>
rect -984 347 984 381
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -381 984 -347
<< locali >>
rect -1180 485 -1084 519
rect 1084 485 1180 519
rect -1180 423 -1146 485
rect 1146 423 1180 485
rect -1000 347 -984 381
rect 984 347 1000 381
rect -1046 297 -1012 313
rect -1046 105 -1012 121
rect 1012 297 1046 313
rect 1012 105 1046 121
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -121 -1012 -105
rect -1046 -313 -1012 -297
rect 1012 -121 1046 -105
rect 1012 -313 1046 -297
rect -1000 -381 -984 -347
rect 984 -381 1000 -347
rect -1180 -485 -1146 -423
rect 1146 -485 1180 -423
rect -1180 -519 -1084 -485
rect 1084 -519 1180 -485
<< viali >>
rect -984 347 984 381
rect -1046 121 -1012 297
rect 1012 121 1046 297
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -297 -1012 -121
rect 1012 -297 1046 -121
rect -984 -381 984 -347
<< metal1 >>
rect -996 381 996 387
rect -996 347 -984 381
rect 984 347 996 381
rect -996 341 996 347
rect -1052 297 -1006 309
rect -1052 121 -1046 297
rect -1012 121 -1006 297
rect -1052 109 -1006 121
rect 1006 297 1052 309
rect 1006 121 1012 297
rect 1046 121 1052 297
rect 1006 109 1052 121
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -121 -1006 -109
rect -1052 -297 -1046 -121
rect -1012 -297 -1006 -121
rect -1052 -309 -1006 -297
rect 1006 -121 1052 -109
rect 1006 -297 1012 -121
rect 1046 -297 1052 -121
rect 1006 -309 1052 -297
rect -996 -347 996 -341
rect -996 -381 -984 -347
rect 984 -381 996 -347
rect -996 -387 996 -381
<< properties >>
string FIXED_BBOX -1163 -502 1163 502
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
