magic
tech sky130A
magscale 1 2
timestamp 1713187236
<< pwell >>
rect -278 -22329 278 22329
<< mvnmos >>
rect -50 20071 50 22071
rect -50 17853 50 19853
rect -50 15635 50 17635
rect -50 13417 50 15417
rect -50 11199 50 13199
rect -50 8981 50 10981
rect -50 6763 50 8763
rect -50 4545 50 6545
rect -50 2327 50 4327
rect -50 109 50 2109
rect -50 -2109 50 -109
rect -50 -4327 50 -2327
rect -50 -6545 50 -4545
rect -50 -8763 50 -6763
rect -50 -10981 50 -8981
rect -50 -13199 50 -11199
rect -50 -15417 50 -13417
rect -50 -17635 50 -15635
rect -50 -19853 50 -17853
rect -50 -22071 50 -20071
<< mvndiff >>
rect -108 22059 -50 22071
rect -108 20083 -96 22059
rect -62 20083 -50 22059
rect -108 20071 -50 20083
rect 50 22059 108 22071
rect 50 20083 62 22059
rect 96 20083 108 22059
rect 50 20071 108 20083
rect -108 19841 -50 19853
rect -108 17865 -96 19841
rect -62 17865 -50 19841
rect -108 17853 -50 17865
rect 50 19841 108 19853
rect 50 17865 62 19841
rect 96 17865 108 19841
rect 50 17853 108 17865
rect -108 17623 -50 17635
rect -108 15647 -96 17623
rect -62 15647 -50 17623
rect -108 15635 -50 15647
rect 50 17623 108 17635
rect 50 15647 62 17623
rect 96 15647 108 17623
rect 50 15635 108 15647
rect -108 15405 -50 15417
rect -108 13429 -96 15405
rect -62 13429 -50 15405
rect -108 13417 -50 13429
rect 50 15405 108 15417
rect 50 13429 62 15405
rect 96 13429 108 15405
rect 50 13417 108 13429
rect -108 13187 -50 13199
rect -108 11211 -96 13187
rect -62 11211 -50 13187
rect -108 11199 -50 11211
rect 50 13187 108 13199
rect 50 11211 62 13187
rect 96 11211 108 13187
rect 50 11199 108 11211
rect -108 10969 -50 10981
rect -108 8993 -96 10969
rect -62 8993 -50 10969
rect -108 8981 -50 8993
rect 50 10969 108 10981
rect 50 8993 62 10969
rect 96 8993 108 10969
rect 50 8981 108 8993
rect -108 8751 -50 8763
rect -108 6775 -96 8751
rect -62 6775 -50 8751
rect -108 6763 -50 6775
rect 50 8751 108 8763
rect 50 6775 62 8751
rect 96 6775 108 8751
rect 50 6763 108 6775
rect -108 6533 -50 6545
rect -108 4557 -96 6533
rect -62 4557 -50 6533
rect -108 4545 -50 4557
rect 50 6533 108 6545
rect 50 4557 62 6533
rect 96 4557 108 6533
rect 50 4545 108 4557
rect -108 4315 -50 4327
rect -108 2339 -96 4315
rect -62 2339 -50 4315
rect -108 2327 -50 2339
rect 50 4315 108 4327
rect 50 2339 62 4315
rect 96 2339 108 4315
rect 50 2327 108 2339
rect -108 2097 -50 2109
rect -108 121 -96 2097
rect -62 121 -50 2097
rect -108 109 -50 121
rect 50 2097 108 2109
rect 50 121 62 2097
rect 96 121 108 2097
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -2097 -96 -121
rect -62 -2097 -50 -121
rect -108 -2109 -50 -2097
rect 50 -121 108 -109
rect 50 -2097 62 -121
rect 96 -2097 108 -121
rect 50 -2109 108 -2097
rect -108 -2339 -50 -2327
rect -108 -4315 -96 -2339
rect -62 -4315 -50 -2339
rect -108 -4327 -50 -4315
rect 50 -2339 108 -2327
rect 50 -4315 62 -2339
rect 96 -4315 108 -2339
rect 50 -4327 108 -4315
rect -108 -4557 -50 -4545
rect -108 -6533 -96 -4557
rect -62 -6533 -50 -4557
rect -108 -6545 -50 -6533
rect 50 -4557 108 -4545
rect 50 -6533 62 -4557
rect 96 -6533 108 -4557
rect 50 -6545 108 -6533
rect -108 -6775 -50 -6763
rect -108 -8751 -96 -6775
rect -62 -8751 -50 -6775
rect -108 -8763 -50 -8751
rect 50 -6775 108 -6763
rect 50 -8751 62 -6775
rect 96 -8751 108 -6775
rect 50 -8763 108 -8751
rect -108 -8993 -50 -8981
rect -108 -10969 -96 -8993
rect -62 -10969 -50 -8993
rect -108 -10981 -50 -10969
rect 50 -8993 108 -8981
rect 50 -10969 62 -8993
rect 96 -10969 108 -8993
rect 50 -10981 108 -10969
rect -108 -11211 -50 -11199
rect -108 -13187 -96 -11211
rect -62 -13187 -50 -11211
rect -108 -13199 -50 -13187
rect 50 -11211 108 -11199
rect 50 -13187 62 -11211
rect 96 -13187 108 -11211
rect 50 -13199 108 -13187
rect -108 -13429 -50 -13417
rect -108 -15405 -96 -13429
rect -62 -15405 -50 -13429
rect -108 -15417 -50 -15405
rect 50 -13429 108 -13417
rect 50 -15405 62 -13429
rect 96 -15405 108 -13429
rect 50 -15417 108 -15405
rect -108 -15647 -50 -15635
rect -108 -17623 -96 -15647
rect -62 -17623 -50 -15647
rect -108 -17635 -50 -17623
rect 50 -15647 108 -15635
rect 50 -17623 62 -15647
rect 96 -17623 108 -15647
rect 50 -17635 108 -17623
rect -108 -17865 -50 -17853
rect -108 -19841 -96 -17865
rect -62 -19841 -50 -17865
rect -108 -19853 -50 -19841
rect 50 -17865 108 -17853
rect 50 -19841 62 -17865
rect 96 -19841 108 -17865
rect 50 -19853 108 -19841
rect -108 -20083 -50 -20071
rect -108 -22059 -96 -20083
rect -62 -22059 -50 -20083
rect -108 -22071 -50 -22059
rect 50 -20083 108 -20071
rect 50 -22059 62 -20083
rect 96 -22059 108 -20083
rect 50 -22071 108 -22059
<< mvndiffc >>
rect -96 20083 -62 22059
rect 62 20083 96 22059
rect -96 17865 -62 19841
rect 62 17865 96 19841
rect -96 15647 -62 17623
rect 62 15647 96 17623
rect -96 13429 -62 15405
rect 62 13429 96 15405
rect -96 11211 -62 13187
rect 62 11211 96 13187
rect -96 8993 -62 10969
rect 62 8993 96 10969
rect -96 6775 -62 8751
rect 62 6775 96 8751
rect -96 4557 -62 6533
rect 62 4557 96 6533
rect -96 2339 -62 4315
rect 62 2339 96 4315
rect -96 121 -62 2097
rect 62 121 96 2097
rect -96 -2097 -62 -121
rect 62 -2097 96 -121
rect -96 -4315 -62 -2339
rect 62 -4315 96 -2339
rect -96 -6533 -62 -4557
rect 62 -6533 96 -4557
rect -96 -8751 -62 -6775
rect 62 -8751 96 -6775
rect -96 -10969 -62 -8993
rect 62 -10969 96 -8993
rect -96 -13187 -62 -11211
rect 62 -13187 96 -11211
rect -96 -15405 -62 -13429
rect 62 -15405 96 -13429
rect -96 -17623 -62 -15647
rect 62 -17623 96 -15647
rect -96 -19841 -62 -17865
rect 62 -19841 96 -17865
rect -96 -22059 -62 -20083
rect 62 -22059 96 -20083
<< mvpsubdiff >>
rect -242 22281 242 22293
rect -242 22247 -134 22281
rect 134 22247 242 22281
rect -242 22235 242 22247
rect -242 22185 -184 22235
rect -242 -22185 -230 22185
rect -196 -22185 -184 22185
rect 184 22185 242 22235
rect -242 -22235 -184 -22185
rect 184 -22185 196 22185
rect 230 -22185 242 22185
rect 184 -22235 242 -22185
rect -242 -22247 242 -22235
rect -242 -22281 -134 -22247
rect 134 -22281 242 -22247
rect -242 -22293 242 -22281
<< mvpsubdiffcont >>
rect -134 22247 134 22281
rect -230 -22185 -196 22185
rect 196 -22185 230 22185
rect -134 -22281 134 -22247
<< poly >>
rect -50 22143 50 22159
rect -50 22109 -34 22143
rect 34 22109 50 22143
rect -50 22071 50 22109
rect -50 20033 50 20071
rect -50 19999 -34 20033
rect 34 19999 50 20033
rect -50 19983 50 19999
rect -50 19925 50 19941
rect -50 19891 -34 19925
rect 34 19891 50 19925
rect -50 19853 50 19891
rect -50 17815 50 17853
rect -50 17781 -34 17815
rect 34 17781 50 17815
rect -50 17765 50 17781
rect -50 17707 50 17723
rect -50 17673 -34 17707
rect 34 17673 50 17707
rect -50 17635 50 17673
rect -50 15597 50 15635
rect -50 15563 -34 15597
rect 34 15563 50 15597
rect -50 15547 50 15563
rect -50 15489 50 15505
rect -50 15455 -34 15489
rect 34 15455 50 15489
rect -50 15417 50 15455
rect -50 13379 50 13417
rect -50 13345 -34 13379
rect 34 13345 50 13379
rect -50 13329 50 13345
rect -50 13271 50 13287
rect -50 13237 -34 13271
rect 34 13237 50 13271
rect -50 13199 50 13237
rect -50 11161 50 11199
rect -50 11127 -34 11161
rect 34 11127 50 11161
rect -50 11111 50 11127
rect -50 11053 50 11069
rect -50 11019 -34 11053
rect 34 11019 50 11053
rect -50 10981 50 11019
rect -50 8943 50 8981
rect -50 8909 -34 8943
rect 34 8909 50 8943
rect -50 8893 50 8909
rect -50 8835 50 8851
rect -50 8801 -34 8835
rect 34 8801 50 8835
rect -50 8763 50 8801
rect -50 6725 50 6763
rect -50 6691 -34 6725
rect 34 6691 50 6725
rect -50 6675 50 6691
rect -50 6617 50 6633
rect -50 6583 -34 6617
rect 34 6583 50 6617
rect -50 6545 50 6583
rect -50 4507 50 4545
rect -50 4473 -34 4507
rect 34 4473 50 4507
rect -50 4457 50 4473
rect -50 4399 50 4415
rect -50 4365 -34 4399
rect 34 4365 50 4399
rect -50 4327 50 4365
rect -50 2289 50 2327
rect -50 2255 -34 2289
rect 34 2255 50 2289
rect -50 2239 50 2255
rect -50 2181 50 2197
rect -50 2147 -34 2181
rect 34 2147 50 2181
rect -50 2109 50 2147
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -2147 50 -2109
rect -50 -2181 -34 -2147
rect 34 -2181 50 -2147
rect -50 -2197 50 -2181
rect -50 -2255 50 -2239
rect -50 -2289 -34 -2255
rect 34 -2289 50 -2255
rect -50 -2327 50 -2289
rect -50 -4365 50 -4327
rect -50 -4399 -34 -4365
rect 34 -4399 50 -4365
rect -50 -4415 50 -4399
rect -50 -4473 50 -4457
rect -50 -4507 -34 -4473
rect 34 -4507 50 -4473
rect -50 -4545 50 -4507
rect -50 -6583 50 -6545
rect -50 -6617 -34 -6583
rect 34 -6617 50 -6583
rect -50 -6633 50 -6617
rect -50 -6691 50 -6675
rect -50 -6725 -34 -6691
rect 34 -6725 50 -6691
rect -50 -6763 50 -6725
rect -50 -8801 50 -8763
rect -50 -8835 -34 -8801
rect 34 -8835 50 -8801
rect -50 -8851 50 -8835
rect -50 -8909 50 -8893
rect -50 -8943 -34 -8909
rect 34 -8943 50 -8909
rect -50 -8981 50 -8943
rect -50 -11019 50 -10981
rect -50 -11053 -34 -11019
rect 34 -11053 50 -11019
rect -50 -11069 50 -11053
rect -50 -11127 50 -11111
rect -50 -11161 -34 -11127
rect 34 -11161 50 -11127
rect -50 -11199 50 -11161
rect -50 -13237 50 -13199
rect -50 -13271 -34 -13237
rect 34 -13271 50 -13237
rect -50 -13287 50 -13271
rect -50 -13345 50 -13329
rect -50 -13379 -34 -13345
rect 34 -13379 50 -13345
rect -50 -13417 50 -13379
rect -50 -15455 50 -15417
rect -50 -15489 -34 -15455
rect 34 -15489 50 -15455
rect -50 -15505 50 -15489
rect -50 -15563 50 -15547
rect -50 -15597 -34 -15563
rect 34 -15597 50 -15563
rect -50 -15635 50 -15597
rect -50 -17673 50 -17635
rect -50 -17707 -34 -17673
rect 34 -17707 50 -17673
rect -50 -17723 50 -17707
rect -50 -17781 50 -17765
rect -50 -17815 -34 -17781
rect 34 -17815 50 -17781
rect -50 -17853 50 -17815
rect -50 -19891 50 -19853
rect -50 -19925 -34 -19891
rect 34 -19925 50 -19891
rect -50 -19941 50 -19925
rect -50 -19999 50 -19983
rect -50 -20033 -34 -19999
rect 34 -20033 50 -19999
rect -50 -20071 50 -20033
rect -50 -22109 50 -22071
rect -50 -22143 -34 -22109
rect 34 -22143 50 -22109
rect -50 -22159 50 -22143
<< polycont >>
rect -34 22109 34 22143
rect -34 19999 34 20033
rect -34 19891 34 19925
rect -34 17781 34 17815
rect -34 17673 34 17707
rect -34 15563 34 15597
rect -34 15455 34 15489
rect -34 13345 34 13379
rect -34 13237 34 13271
rect -34 11127 34 11161
rect -34 11019 34 11053
rect -34 8909 34 8943
rect -34 8801 34 8835
rect -34 6691 34 6725
rect -34 6583 34 6617
rect -34 4473 34 4507
rect -34 4365 34 4399
rect -34 2255 34 2289
rect -34 2147 34 2181
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -2181 34 -2147
rect -34 -2289 34 -2255
rect -34 -4399 34 -4365
rect -34 -4507 34 -4473
rect -34 -6617 34 -6583
rect -34 -6725 34 -6691
rect -34 -8835 34 -8801
rect -34 -8943 34 -8909
rect -34 -11053 34 -11019
rect -34 -11161 34 -11127
rect -34 -13271 34 -13237
rect -34 -13379 34 -13345
rect -34 -15489 34 -15455
rect -34 -15597 34 -15563
rect -34 -17707 34 -17673
rect -34 -17815 34 -17781
rect -34 -19925 34 -19891
rect -34 -20033 34 -19999
rect -34 -22143 34 -22109
<< locali >>
rect -230 22247 -134 22281
rect 134 22247 230 22281
rect -230 22185 -196 22247
rect 196 22185 230 22247
rect -50 22109 -34 22143
rect 34 22109 50 22143
rect -96 22059 -62 22075
rect -96 20067 -62 20083
rect 62 22059 96 22075
rect 62 20067 96 20083
rect -50 19999 -34 20033
rect 34 19999 50 20033
rect -50 19891 -34 19925
rect 34 19891 50 19925
rect -96 19841 -62 19857
rect -96 17849 -62 17865
rect 62 19841 96 19857
rect 62 17849 96 17865
rect -50 17781 -34 17815
rect 34 17781 50 17815
rect -50 17673 -34 17707
rect 34 17673 50 17707
rect -96 17623 -62 17639
rect -96 15631 -62 15647
rect 62 17623 96 17639
rect 62 15631 96 15647
rect -50 15563 -34 15597
rect 34 15563 50 15597
rect -50 15455 -34 15489
rect 34 15455 50 15489
rect -96 15405 -62 15421
rect -96 13413 -62 13429
rect 62 15405 96 15421
rect 62 13413 96 13429
rect -50 13345 -34 13379
rect 34 13345 50 13379
rect -50 13237 -34 13271
rect 34 13237 50 13271
rect -96 13187 -62 13203
rect -96 11195 -62 11211
rect 62 13187 96 13203
rect 62 11195 96 11211
rect -50 11127 -34 11161
rect 34 11127 50 11161
rect -50 11019 -34 11053
rect 34 11019 50 11053
rect -96 10969 -62 10985
rect -96 8977 -62 8993
rect 62 10969 96 10985
rect 62 8977 96 8993
rect -50 8909 -34 8943
rect 34 8909 50 8943
rect -50 8801 -34 8835
rect 34 8801 50 8835
rect -96 8751 -62 8767
rect -96 6759 -62 6775
rect 62 8751 96 8767
rect 62 6759 96 6775
rect -50 6691 -34 6725
rect 34 6691 50 6725
rect -50 6583 -34 6617
rect 34 6583 50 6617
rect -96 6533 -62 6549
rect -96 4541 -62 4557
rect 62 6533 96 6549
rect 62 4541 96 4557
rect -50 4473 -34 4507
rect 34 4473 50 4507
rect -50 4365 -34 4399
rect 34 4365 50 4399
rect -96 4315 -62 4331
rect -96 2323 -62 2339
rect 62 4315 96 4331
rect 62 2323 96 2339
rect -50 2255 -34 2289
rect 34 2255 50 2289
rect -50 2147 -34 2181
rect 34 2147 50 2181
rect -96 2097 -62 2113
rect -96 105 -62 121
rect 62 2097 96 2113
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -2113 -62 -2097
rect 62 -121 96 -105
rect 62 -2113 96 -2097
rect -50 -2181 -34 -2147
rect 34 -2181 50 -2147
rect -50 -2289 -34 -2255
rect 34 -2289 50 -2255
rect -96 -2339 -62 -2323
rect -96 -4331 -62 -4315
rect 62 -2339 96 -2323
rect 62 -4331 96 -4315
rect -50 -4399 -34 -4365
rect 34 -4399 50 -4365
rect -50 -4507 -34 -4473
rect 34 -4507 50 -4473
rect -96 -4557 -62 -4541
rect -96 -6549 -62 -6533
rect 62 -4557 96 -4541
rect 62 -6549 96 -6533
rect -50 -6617 -34 -6583
rect 34 -6617 50 -6583
rect -50 -6725 -34 -6691
rect 34 -6725 50 -6691
rect -96 -6775 -62 -6759
rect -96 -8767 -62 -8751
rect 62 -6775 96 -6759
rect 62 -8767 96 -8751
rect -50 -8835 -34 -8801
rect 34 -8835 50 -8801
rect -50 -8943 -34 -8909
rect 34 -8943 50 -8909
rect -96 -8993 -62 -8977
rect -96 -10985 -62 -10969
rect 62 -8993 96 -8977
rect 62 -10985 96 -10969
rect -50 -11053 -34 -11019
rect 34 -11053 50 -11019
rect -50 -11161 -34 -11127
rect 34 -11161 50 -11127
rect -96 -11211 -62 -11195
rect -96 -13203 -62 -13187
rect 62 -11211 96 -11195
rect 62 -13203 96 -13187
rect -50 -13271 -34 -13237
rect 34 -13271 50 -13237
rect -50 -13379 -34 -13345
rect 34 -13379 50 -13345
rect -96 -13429 -62 -13413
rect -96 -15421 -62 -15405
rect 62 -13429 96 -13413
rect 62 -15421 96 -15405
rect -50 -15489 -34 -15455
rect 34 -15489 50 -15455
rect -50 -15597 -34 -15563
rect 34 -15597 50 -15563
rect -96 -15647 -62 -15631
rect -96 -17639 -62 -17623
rect 62 -15647 96 -15631
rect 62 -17639 96 -17623
rect -50 -17707 -34 -17673
rect 34 -17707 50 -17673
rect -50 -17815 -34 -17781
rect 34 -17815 50 -17781
rect -96 -17865 -62 -17849
rect -96 -19857 -62 -19841
rect 62 -17865 96 -17849
rect 62 -19857 96 -19841
rect -50 -19925 -34 -19891
rect 34 -19925 50 -19891
rect -50 -20033 -34 -19999
rect 34 -20033 50 -19999
rect -96 -20083 -62 -20067
rect -96 -22075 -62 -22059
rect 62 -20083 96 -20067
rect 62 -22075 96 -22059
rect -50 -22143 -34 -22109
rect 34 -22143 50 -22109
rect -230 -22247 -196 -22185
rect 196 -22247 230 -22185
rect -230 -22281 -134 -22247
rect 134 -22281 230 -22247
<< viali >>
rect -34 22109 34 22143
rect -96 20083 -62 22059
rect 62 20083 96 22059
rect -34 19999 34 20033
rect -34 19891 34 19925
rect -96 17865 -62 19841
rect 62 17865 96 19841
rect -34 17781 34 17815
rect -34 17673 34 17707
rect -96 15647 -62 17623
rect 62 15647 96 17623
rect -34 15563 34 15597
rect -34 15455 34 15489
rect -96 13429 -62 15405
rect 62 13429 96 15405
rect -34 13345 34 13379
rect -34 13237 34 13271
rect -96 11211 -62 13187
rect 62 11211 96 13187
rect -34 11127 34 11161
rect -34 11019 34 11053
rect -96 8993 -62 10969
rect 62 8993 96 10969
rect -34 8909 34 8943
rect -34 8801 34 8835
rect -96 6775 -62 8751
rect 62 6775 96 8751
rect -34 6691 34 6725
rect -34 6583 34 6617
rect -96 4557 -62 6533
rect 62 4557 96 6533
rect -34 4473 34 4507
rect -34 4365 34 4399
rect -96 2339 -62 4315
rect 62 2339 96 4315
rect -34 2255 34 2289
rect -34 2147 34 2181
rect -96 121 -62 2097
rect 62 121 96 2097
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -2097 -62 -121
rect 62 -2097 96 -121
rect -34 -2181 34 -2147
rect -34 -2289 34 -2255
rect -96 -4315 -62 -2339
rect 62 -4315 96 -2339
rect -34 -4399 34 -4365
rect -34 -4507 34 -4473
rect -96 -6533 -62 -4557
rect 62 -6533 96 -4557
rect -34 -6617 34 -6583
rect -34 -6725 34 -6691
rect -96 -8751 -62 -6775
rect 62 -8751 96 -6775
rect -34 -8835 34 -8801
rect -34 -8943 34 -8909
rect -96 -10969 -62 -8993
rect 62 -10969 96 -8993
rect -34 -11053 34 -11019
rect -34 -11161 34 -11127
rect -96 -13187 -62 -11211
rect 62 -13187 96 -11211
rect -34 -13271 34 -13237
rect -34 -13379 34 -13345
rect -96 -15405 -62 -13429
rect 62 -15405 96 -13429
rect -34 -15489 34 -15455
rect -34 -15597 34 -15563
rect -96 -17623 -62 -15647
rect 62 -17623 96 -15647
rect -34 -17707 34 -17673
rect -34 -17815 34 -17781
rect -96 -19841 -62 -17865
rect 62 -19841 96 -17865
rect -34 -19925 34 -19891
rect -34 -20033 34 -19999
rect -96 -22059 -62 -20083
rect 62 -22059 96 -20083
rect -34 -22143 34 -22109
<< metal1 >>
rect -46 22143 46 22149
rect -46 22109 -34 22143
rect 34 22109 46 22143
rect -46 22103 46 22109
rect -102 22059 -56 22071
rect -102 20083 -96 22059
rect -62 20083 -56 22059
rect -102 20071 -56 20083
rect 56 22059 102 22071
rect 56 20083 62 22059
rect 96 20083 102 22059
rect 56 20071 102 20083
rect -46 20033 46 20039
rect -46 19999 -34 20033
rect 34 19999 46 20033
rect -46 19993 46 19999
rect -46 19925 46 19931
rect -46 19891 -34 19925
rect 34 19891 46 19925
rect -46 19885 46 19891
rect -102 19841 -56 19853
rect -102 17865 -96 19841
rect -62 17865 -56 19841
rect -102 17853 -56 17865
rect 56 19841 102 19853
rect 56 17865 62 19841
rect 96 17865 102 19841
rect 56 17853 102 17865
rect -46 17815 46 17821
rect -46 17781 -34 17815
rect 34 17781 46 17815
rect -46 17775 46 17781
rect -46 17707 46 17713
rect -46 17673 -34 17707
rect 34 17673 46 17707
rect -46 17667 46 17673
rect -102 17623 -56 17635
rect -102 15647 -96 17623
rect -62 15647 -56 17623
rect -102 15635 -56 15647
rect 56 17623 102 17635
rect 56 15647 62 17623
rect 96 15647 102 17623
rect 56 15635 102 15647
rect -46 15597 46 15603
rect -46 15563 -34 15597
rect 34 15563 46 15597
rect -46 15557 46 15563
rect -46 15489 46 15495
rect -46 15455 -34 15489
rect 34 15455 46 15489
rect -46 15449 46 15455
rect -102 15405 -56 15417
rect -102 13429 -96 15405
rect -62 13429 -56 15405
rect -102 13417 -56 13429
rect 56 15405 102 15417
rect 56 13429 62 15405
rect 96 13429 102 15405
rect 56 13417 102 13429
rect -46 13379 46 13385
rect -46 13345 -34 13379
rect 34 13345 46 13379
rect -46 13339 46 13345
rect -46 13271 46 13277
rect -46 13237 -34 13271
rect 34 13237 46 13271
rect -46 13231 46 13237
rect -102 13187 -56 13199
rect -102 11211 -96 13187
rect -62 11211 -56 13187
rect -102 11199 -56 11211
rect 56 13187 102 13199
rect 56 11211 62 13187
rect 96 11211 102 13187
rect 56 11199 102 11211
rect -46 11161 46 11167
rect -46 11127 -34 11161
rect 34 11127 46 11161
rect -46 11121 46 11127
rect -46 11053 46 11059
rect -46 11019 -34 11053
rect 34 11019 46 11053
rect -46 11013 46 11019
rect -102 10969 -56 10981
rect -102 8993 -96 10969
rect -62 8993 -56 10969
rect -102 8981 -56 8993
rect 56 10969 102 10981
rect 56 8993 62 10969
rect 96 8993 102 10969
rect 56 8981 102 8993
rect -46 8943 46 8949
rect -46 8909 -34 8943
rect 34 8909 46 8943
rect -46 8903 46 8909
rect -46 8835 46 8841
rect -46 8801 -34 8835
rect 34 8801 46 8835
rect -46 8795 46 8801
rect -102 8751 -56 8763
rect -102 6775 -96 8751
rect -62 6775 -56 8751
rect -102 6763 -56 6775
rect 56 8751 102 8763
rect 56 6775 62 8751
rect 96 6775 102 8751
rect 56 6763 102 6775
rect -46 6725 46 6731
rect -46 6691 -34 6725
rect 34 6691 46 6725
rect -46 6685 46 6691
rect -46 6617 46 6623
rect -46 6583 -34 6617
rect 34 6583 46 6617
rect -46 6577 46 6583
rect -102 6533 -56 6545
rect -102 4557 -96 6533
rect -62 4557 -56 6533
rect -102 4545 -56 4557
rect 56 6533 102 6545
rect 56 4557 62 6533
rect 96 4557 102 6533
rect 56 4545 102 4557
rect -46 4507 46 4513
rect -46 4473 -34 4507
rect 34 4473 46 4507
rect -46 4467 46 4473
rect -46 4399 46 4405
rect -46 4365 -34 4399
rect 34 4365 46 4399
rect -46 4359 46 4365
rect -102 4315 -56 4327
rect -102 2339 -96 4315
rect -62 2339 -56 4315
rect -102 2327 -56 2339
rect 56 4315 102 4327
rect 56 2339 62 4315
rect 96 2339 102 4315
rect 56 2327 102 2339
rect -46 2289 46 2295
rect -46 2255 -34 2289
rect 34 2255 46 2289
rect -46 2249 46 2255
rect -46 2181 46 2187
rect -46 2147 -34 2181
rect 34 2147 46 2181
rect -46 2141 46 2147
rect -102 2097 -56 2109
rect -102 121 -96 2097
rect -62 121 -56 2097
rect -102 109 -56 121
rect 56 2097 102 2109
rect 56 121 62 2097
rect 96 121 102 2097
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -2097 -96 -121
rect -62 -2097 -56 -121
rect -102 -2109 -56 -2097
rect 56 -121 102 -109
rect 56 -2097 62 -121
rect 96 -2097 102 -121
rect 56 -2109 102 -2097
rect -46 -2147 46 -2141
rect -46 -2181 -34 -2147
rect 34 -2181 46 -2147
rect -46 -2187 46 -2181
rect -46 -2255 46 -2249
rect -46 -2289 -34 -2255
rect 34 -2289 46 -2255
rect -46 -2295 46 -2289
rect -102 -2339 -56 -2327
rect -102 -4315 -96 -2339
rect -62 -4315 -56 -2339
rect -102 -4327 -56 -4315
rect 56 -2339 102 -2327
rect 56 -4315 62 -2339
rect 96 -4315 102 -2339
rect 56 -4327 102 -4315
rect -46 -4365 46 -4359
rect -46 -4399 -34 -4365
rect 34 -4399 46 -4365
rect -46 -4405 46 -4399
rect -46 -4473 46 -4467
rect -46 -4507 -34 -4473
rect 34 -4507 46 -4473
rect -46 -4513 46 -4507
rect -102 -4557 -56 -4545
rect -102 -6533 -96 -4557
rect -62 -6533 -56 -4557
rect -102 -6545 -56 -6533
rect 56 -4557 102 -4545
rect 56 -6533 62 -4557
rect 96 -6533 102 -4557
rect 56 -6545 102 -6533
rect -46 -6583 46 -6577
rect -46 -6617 -34 -6583
rect 34 -6617 46 -6583
rect -46 -6623 46 -6617
rect -46 -6691 46 -6685
rect -46 -6725 -34 -6691
rect 34 -6725 46 -6691
rect -46 -6731 46 -6725
rect -102 -6775 -56 -6763
rect -102 -8751 -96 -6775
rect -62 -8751 -56 -6775
rect -102 -8763 -56 -8751
rect 56 -6775 102 -6763
rect 56 -8751 62 -6775
rect 96 -8751 102 -6775
rect 56 -8763 102 -8751
rect -46 -8801 46 -8795
rect -46 -8835 -34 -8801
rect 34 -8835 46 -8801
rect -46 -8841 46 -8835
rect -46 -8909 46 -8903
rect -46 -8943 -34 -8909
rect 34 -8943 46 -8909
rect -46 -8949 46 -8943
rect -102 -8993 -56 -8981
rect -102 -10969 -96 -8993
rect -62 -10969 -56 -8993
rect -102 -10981 -56 -10969
rect 56 -8993 102 -8981
rect 56 -10969 62 -8993
rect 96 -10969 102 -8993
rect 56 -10981 102 -10969
rect -46 -11019 46 -11013
rect -46 -11053 -34 -11019
rect 34 -11053 46 -11019
rect -46 -11059 46 -11053
rect -46 -11127 46 -11121
rect -46 -11161 -34 -11127
rect 34 -11161 46 -11127
rect -46 -11167 46 -11161
rect -102 -11211 -56 -11199
rect -102 -13187 -96 -11211
rect -62 -13187 -56 -11211
rect -102 -13199 -56 -13187
rect 56 -11211 102 -11199
rect 56 -13187 62 -11211
rect 96 -13187 102 -11211
rect 56 -13199 102 -13187
rect -46 -13237 46 -13231
rect -46 -13271 -34 -13237
rect 34 -13271 46 -13237
rect -46 -13277 46 -13271
rect -46 -13345 46 -13339
rect -46 -13379 -34 -13345
rect 34 -13379 46 -13345
rect -46 -13385 46 -13379
rect -102 -13429 -56 -13417
rect -102 -15405 -96 -13429
rect -62 -15405 -56 -13429
rect -102 -15417 -56 -15405
rect 56 -13429 102 -13417
rect 56 -15405 62 -13429
rect 96 -15405 102 -13429
rect 56 -15417 102 -15405
rect -46 -15455 46 -15449
rect -46 -15489 -34 -15455
rect 34 -15489 46 -15455
rect -46 -15495 46 -15489
rect -46 -15563 46 -15557
rect -46 -15597 -34 -15563
rect 34 -15597 46 -15563
rect -46 -15603 46 -15597
rect -102 -15647 -56 -15635
rect -102 -17623 -96 -15647
rect -62 -17623 -56 -15647
rect -102 -17635 -56 -17623
rect 56 -15647 102 -15635
rect 56 -17623 62 -15647
rect 96 -17623 102 -15647
rect 56 -17635 102 -17623
rect -46 -17673 46 -17667
rect -46 -17707 -34 -17673
rect 34 -17707 46 -17673
rect -46 -17713 46 -17707
rect -46 -17781 46 -17775
rect -46 -17815 -34 -17781
rect 34 -17815 46 -17781
rect -46 -17821 46 -17815
rect -102 -17865 -56 -17853
rect -102 -19841 -96 -17865
rect -62 -19841 -56 -17865
rect -102 -19853 -56 -19841
rect 56 -17865 102 -17853
rect 56 -19841 62 -17865
rect 96 -19841 102 -17865
rect 56 -19853 102 -19841
rect -46 -19891 46 -19885
rect -46 -19925 -34 -19891
rect 34 -19925 46 -19891
rect -46 -19931 46 -19925
rect -46 -19999 46 -19993
rect -46 -20033 -34 -19999
rect 34 -20033 46 -19999
rect -46 -20039 46 -20033
rect -102 -20083 -56 -20071
rect -102 -22059 -96 -20083
rect -62 -22059 -56 -20083
rect -102 -22071 -56 -22059
rect 56 -20083 102 -20071
rect 56 -22059 62 -20083
rect 96 -22059 102 -20083
rect 56 -22071 102 -22059
rect -46 -22109 46 -22103
rect -46 -22143 -34 -22109
rect 34 -22143 46 -22109
rect -46 -22149 46 -22143
<< properties >>
string FIXED_BBOX -213 -22264 213 22264
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
