magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -1258 -1487 1258 1487
<< mvpmos >>
rect -1000 990 1000 1190
rect -1000 554 1000 754
rect -1000 118 1000 318
rect -1000 -318 1000 -118
rect -1000 -754 1000 -554
rect -1000 -1190 1000 -990
<< mvpdiff >>
rect -1058 1178 -1000 1190
rect -1058 1002 -1046 1178
rect -1012 1002 -1000 1178
rect -1058 990 -1000 1002
rect 1000 1178 1058 1190
rect 1000 1002 1012 1178
rect 1046 1002 1058 1178
rect 1000 990 1058 1002
rect -1058 742 -1000 754
rect -1058 566 -1046 742
rect -1012 566 -1000 742
rect -1058 554 -1000 566
rect 1000 742 1058 754
rect 1000 566 1012 742
rect 1046 566 1058 742
rect 1000 554 1058 566
rect -1058 306 -1000 318
rect -1058 130 -1046 306
rect -1012 130 -1000 306
rect -1058 118 -1000 130
rect 1000 306 1058 318
rect 1000 130 1012 306
rect 1046 130 1058 306
rect 1000 118 1058 130
rect -1058 -130 -1000 -118
rect -1058 -306 -1046 -130
rect -1012 -306 -1000 -130
rect -1058 -318 -1000 -306
rect 1000 -130 1058 -118
rect 1000 -306 1012 -130
rect 1046 -306 1058 -130
rect 1000 -318 1058 -306
rect -1058 -566 -1000 -554
rect -1058 -742 -1046 -566
rect -1012 -742 -1000 -566
rect -1058 -754 -1000 -742
rect 1000 -566 1058 -554
rect 1000 -742 1012 -566
rect 1046 -742 1058 -566
rect 1000 -754 1058 -742
rect -1058 -1002 -1000 -990
rect -1058 -1178 -1046 -1002
rect -1012 -1178 -1000 -1002
rect -1058 -1190 -1000 -1178
rect 1000 -1002 1058 -990
rect 1000 -1178 1012 -1002
rect 1046 -1178 1058 -1002
rect 1000 -1190 1058 -1178
<< mvpdiffc >>
rect -1046 1002 -1012 1178
rect 1012 1002 1046 1178
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
rect -1046 -1178 -1012 -1002
rect 1012 -1178 1046 -1002
<< mvnsubdiff >>
rect -1192 1409 1192 1421
rect -1192 1375 -1084 1409
rect 1084 1375 1192 1409
rect -1192 1363 1192 1375
rect -1192 1313 -1134 1363
rect -1192 -1313 -1180 1313
rect -1146 -1313 -1134 1313
rect 1134 1313 1192 1363
rect -1192 -1363 -1134 -1313
rect 1134 -1313 1146 1313
rect 1180 -1313 1192 1313
rect 1134 -1363 1192 -1313
rect -1192 -1375 1192 -1363
rect -1192 -1409 -1084 -1375
rect 1084 -1409 1192 -1375
rect -1192 -1421 1192 -1409
<< mvnsubdiffcont >>
rect -1084 1375 1084 1409
rect -1180 -1313 -1146 1313
rect 1146 -1313 1180 1313
rect -1084 -1409 1084 -1375
<< poly >>
rect -1000 1271 1000 1287
rect -1000 1237 -984 1271
rect 984 1237 1000 1271
rect -1000 1190 1000 1237
rect -1000 943 1000 990
rect -1000 909 -984 943
rect 984 909 1000 943
rect -1000 893 1000 909
rect -1000 835 1000 851
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1000 754 1000 801
rect -1000 507 1000 554
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 457 1000 473
rect -1000 399 1000 415
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1000 318 1000 365
rect -1000 71 1000 118
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -118 1000 -71
rect -1000 -365 1000 -318
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -415 1000 -399
rect -1000 -473 1000 -457
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1000 -554 1000 -507
rect -1000 -801 1000 -754
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect -1000 -851 1000 -835
rect -1000 -909 1000 -893
rect -1000 -943 -984 -909
rect 984 -943 1000 -909
rect -1000 -990 1000 -943
rect -1000 -1237 1000 -1190
rect -1000 -1271 -984 -1237
rect 984 -1271 1000 -1237
rect -1000 -1287 1000 -1271
<< polycont >>
rect -984 1237 984 1271
rect -984 909 984 943
rect -984 801 984 835
rect -984 473 984 507
rect -984 365 984 399
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -399 984 -365
rect -984 -507 984 -473
rect -984 -835 984 -801
rect -984 -943 984 -909
rect -984 -1271 984 -1237
<< locali >>
rect -1180 1375 -1084 1409
rect 1084 1375 1180 1409
rect -1180 1313 -1146 1375
rect 1146 1313 1180 1375
rect -1000 1237 -984 1271
rect 984 1237 1000 1271
rect -1046 1178 -1012 1194
rect -1046 986 -1012 1002
rect 1012 1178 1046 1194
rect 1012 986 1046 1002
rect -1000 909 -984 943
rect 984 909 1000 943
rect -1000 801 -984 835
rect 984 801 1000 835
rect -1046 742 -1012 758
rect -1046 550 -1012 566
rect 1012 742 1046 758
rect 1012 550 1046 566
rect -1000 473 -984 507
rect 984 473 1000 507
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1046 306 -1012 322
rect -1046 114 -1012 130
rect 1012 306 1046 322
rect 1012 114 1046 130
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -130 -1012 -114
rect -1046 -322 -1012 -306
rect 1012 -130 1046 -114
rect 1012 -322 1046 -306
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -507 -984 -473
rect 984 -507 1000 -473
rect -1046 -566 -1012 -550
rect -1046 -758 -1012 -742
rect 1012 -566 1046 -550
rect 1012 -758 1046 -742
rect -1000 -835 -984 -801
rect 984 -835 1000 -801
rect -1000 -943 -984 -909
rect 984 -943 1000 -909
rect -1046 -1002 -1012 -986
rect -1046 -1194 -1012 -1178
rect 1012 -1002 1046 -986
rect 1012 -1194 1046 -1178
rect -1000 -1271 -984 -1237
rect 984 -1271 1000 -1237
rect -1180 -1375 -1146 -1313
rect 1146 -1375 1180 -1313
rect -1180 -1409 -1084 -1375
rect 1084 -1409 1180 -1375
<< viali >>
rect -984 1237 984 1271
rect -1046 1002 -1012 1178
rect 1012 1002 1046 1178
rect -984 909 984 943
rect -984 801 984 835
rect -1046 566 -1012 742
rect 1012 566 1046 742
rect -984 473 984 507
rect -984 365 984 399
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -984 -399 984 -365
rect -984 -507 984 -473
rect -1046 -742 -1012 -566
rect 1012 -742 1046 -566
rect -984 -835 984 -801
rect -984 -943 984 -909
rect -1046 -1178 -1012 -1002
rect 1012 -1178 1046 -1002
rect -984 -1271 984 -1237
<< metal1 >>
rect -996 1271 996 1277
rect -996 1237 -984 1271
rect 984 1237 996 1271
rect -996 1231 996 1237
rect -1052 1178 -1006 1190
rect -1052 1002 -1046 1178
rect -1012 1002 -1006 1178
rect -1052 990 -1006 1002
rect 1006 1178 1052 1190
rect 1006 1002 1012 1178
rect 1046 1002 1052 1178
rect 1006 990 1052 1002
rect -996 943 996 949
rect -996 909 -984 943
rect 984 909 996 943
rect -996 903 996 909
rect -996 835 996 841
rect -996 801 -984 835
rect 984 801 996 835
rect -996 795 996 801
rect -1052 742 -1006 754
rect -1052 566 -1046 742
rect -1012 566 -1006 742
rect -1052 554 -1006 566
rect 1006 742 1052 754
rect 1006 566 1012 742
rect 1046 566 1052 742
rect 1006 554 1052 566
rect -996 507 996 513
rect -996 473 -984 507
rect 984 473 996 507
rect -996 467 996 473
rect -996 399 996 405
rect -996 365 -984 399
rect 984 365 996 399
rect -996 359 996 365
rect -1052 306 -1006 318
rect -1052 130 -1046 306
rect -1012 130 -1006 306
rect -1052 118 -1006 130
rect 1006 306 1052 318
rect 1006 130 1012 306
rect 1046 130 1052 306
rect 1006 118 1052 130
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -130 -1006 -118
rect -1052 -306 -1046 -130
rect -1012 -306 -1006 -130
rect -1052 -318 -1006 -306
rect 1006 -130 1052 -118
rect 1006 -306 1012 -130
rect 1046 -306 1052 -130
rect 1006 -318 1052 -306
rect -996 -365 996 -359
rect -996 -399 -984 -365
rect 984 -399 996 -365
rect -996 -405 996 -399
rect -996 -473 996 -467
rect -996 -507 -984 -473
rect 984 -507 996 -473
rect -996 -513 996 -507
rect -1052 -566 -1006 -554
rect -1052 -742 -1046 -566
rect -1012 -742 -1006 -566
rect -1052 -754 -1006 -742
rect 1006 -566 1052 -554
rect 1006 -742 1012 -566
rect 1046 -742 1052 -566
rect 1006 -754 1052 -742
rect -996 -801 996 -795
rect -996 -835 -984 -801
rect 984 -835 996 -801
rect -996 -841 996 -835
rect -996 -909 996 -903
rect -996 -943 -984 -909
rect 984 -943 996 -909
rect -996 -949 996 -943
rect -1052 -1002 -1006 -990
rect -1052 -1178 -1046 -1002
rect -1012 -1178 -1006 -1002
rect -1052 -1190 -1006 -1178
rect 1006 -1002 1052 -990
rect 1006 -1178 1012 -1002
rect 1046 -1178 1052 -1002
rect 1006 -1190 1052 -1178
rect -996 -1237 996 -1231
rect -996 -1271 -984 -1237
rect 984 -1271 996 -1237
rect -996 -1277 996 -1271
<< properties >>
string FIXED_BBOX -1163 -1392 1163 1392
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
