magic
tech sky130A
magscale 1 2
timestamp 1717253844
<< pwell >>
rect -201 -36582 201 36582
<< psubdiff >>
rect -165 36512 -69 36546
rect 69 36512 165 36546
rect -165 36450 -131 36512
rect 131 36450 165 36512
rect -165 -36512 -131 -36450
rect 131 -36512 165 -36450
rect -165 -36546 -69 -36512
rect 69 -36546 165 -36512
<< psubdiffcont >>
rect -69 36512 69 36546
rect -165 -36450 -131 36450
rect 131 -36450 165 36450
rect -69 -36546 69 -36512
<< xpolycontact >>
rect -35 35984 35 36416
rect -35 -36416 35 -35984
<< xpolyres >>
rect -35 -35984 35 35984
<< locali >>
rect -165 36512 -69 36546
rect 69 36512 165 36546
rect -165 36450 -131 36512
rect 131 36450 165 36512
rect -165 -36512 -131 -36450
rect 131 -36512 165 -36450
rect -165 -36546 -69 -36512
rect 69 -36546 165 -36512
<< viali >>
rect -19 36001 19 36398
rect -19 -36398 19 -36001
<< metal1 >>
rect -25 36398 25 36410
rect -25 36001 -19 36398
rect 19 36001 25 36398
rect -25 35989 25 36001
rect -25 -36001 25 -35989
rect -25 -36398 -19 -36001
rect 19 -36398 25 -36001
rect -25 -36410 25 -36398
<< properties >>
string FIXED_BBOX -148 -36529 148 36529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 360.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 2.058meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
