magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -1258 -3449 1258 3449
<< mvpmos >>
rect -1000 2952 1000 3152
rect -1000 2516 1000 2716
rect -1000 2080 1000 2280
rect -1000 1644 1000 1844
rect -1000 1208 1000 1408
rect -1000 772 1000 972
rect -1000 336 1000 536
rect -1000 -100 1000 100
rect -1000 -536 1000 -336
rect -1000 -972 1000 -772
rect -1000 -1408 1000 -1208
rect -1000 -1844 1000 -1644
rect -1000 -2280 1000 -2080
rect -1000 -2716 1000 -2516
rect -1000 -3152 1000 -2952
<< mvpdiff >>
rect -1058 3140 -1000 3152
rect -1058 2964 -1046 3140
rect -1012 2964 -1000 3140
rect -1058 2952 -1000 2964
rect 1000 3140 1058 3152
rect 1000 2964 1012 3140
rect 1046 2964 1058 3140
rect 1000 2952 1058 2964
rect -1058 2704 -1000 2716
rect -1058 2528 -1046 2704
rect -1012 2528 -1000 2704
rect -1058 2516 -1000 2528
rect 1000 2704 1058 2716
rect 1000 2528 1012 2704
rect 1046 2528 1058 2704
rect 1000 2516 1058 2528
rect -1058 2268 -1000 2280
rect -1058 2092 -1046 2268
rect -1012 2092 -1000 2268
rect -1058 2080 -1000 2092
rect 1000 2268 1058 2280
rect 1000 2092 1012 2268
rect 1046 2092 1058 2268
rect 1000 2080 1058 2092
rect -1058 1832 -1000 1844
rect -1058 1656 -1046 1832
rect -1012 1656 -1000 1832
rect -1058 1644 -1000 1656
rect 1000 1832 1058 1844
rect 1000 1656 1012 1832
rect 1046 1656 1058 1832
rect 1000 1644 1058 1656
rect -1058 1396 -1000 1408
rect -1058 1220 -1046 1396
rect -1012 1220 -1000 1396
rect -1058 1208 -1000 1220
rect 1000 1396 1058 1408
rect 1000 1220 1012 1396
rect 1046 1220 1058 1396
rect 1000 1208 1058 1220
rect -1058 960 -1000 972
rect -1058 784 -1046 960
rect -1012 784 -1000 960
rect -1058 772 -1000 784
rect 1000 960 1058 972
rect 1000 784 1012 960
rect 1046 784 1058 960
rect 1000 772 1058 784
rect -1058 524 -1000 536
rect -1058 348 -1046 524
rect -1012 348 -1000 524
rect -1058 336 -1000 348
rect 1000 524 1058 536
rect 1000 348 1012 524
rect 1046 348 1058 524
rect 1000 336 1058 348
rect -1058 88 -1000 100
rect -1058 -88 -1046 88
rect -1012 -88 -1000 88
rect -1058 -100 -1000 -88
rect 1000 88 1058 100
rect 1000 -88 1012 88
rect 1046 -88 1058 88
rect 1000 -100 1058 -88
rect -1058 -348 -1000 -336
rect -1058 -524 -1046 -348
rect -1012 -524 -1000 -348
rect -1058 -536 -1000 -524
rect 1000 -348 1058 -336
rect 1000 -524 1012 -348
rect 1046 -524 1058 -348
rect 1000 -536 1058 -524
rect -1058 -784 -1000 -772
rect -1058 -960 -1046 -784
rect -1012 -960 -1000 -784
rect -1058 -972 -1000 -960
rect 1000 -784 1058 -772
rect 1000 -960 1012 -784
rect 1046 -960 1058 -784
rect 1000 -972 1058 -960
rect -1058 -1220 -1000 -1208
rect -1058 -1396 -1046 -1220
rect -1012 -1396 -1000 -1220
rect -1058 -1408 -1000 -1396
rect 1000 -1220 1058 -1208
rect 1000 -1396 1012 -1220
rect 1046 -1396 1058 -1220
rect 1000 -1408 1058 -1396
rect -1058 -1656 -1000 -1644
rect -1058 -1832 -1046 -1656
rect -1012 -1832 -1000 -1656
rect -1058 -1844 -1000 -1832
rect 1000 -1656 1058 -1644
rect 1000 -1832 1012 -1656
rect 1046 -1832 1058 -1656
rect 1000 -1844 1058 -1832
rect -1058 -2092 -1000 -2080
rect -1058 -2268 -1046 -2092
rect -1012 -2268 -1000 -2092
rect -1058 -2280 -1000 -2268
rect 1000 -2092 1058 -2080
rect 1000 -2268 1012 -2092
rect 1046 -2268 1058 -2092
rect 1000 -2280 1058 -2268
rect -1058 -2528 -1000 -2516
rect -1058 -2704 -1046 -2528
rect -1012 -2704 -1000 -2528
rect -1058 -2716 -1000 -2704
rect 1000 -2528 1058 -2516
rect 1000 -2704 1012 -2528
rect 1046 -2704 1058 -2528
rect 1000 -2716 1058 -2704
rect -1058 -2964 -1000 -2952
rect -1058 -3140 -1046 -2964
rect -1012 -3140 -1000 -2964
rect -1058 -3152 -1000 -3140
rect 1000 -2964 1058 -2952
rect 1000 -3140 1012 -2964
rect 1046 -3140 1058 -2964
rect 1000 -3152 1058 -3140
<< mvpdiffc >>
rect -1046 2964 -1012 3140
rect 1012 2964 1046 3140
rect -1046 2528 -1012 2704
rect 1012 2528 1046 2704
rect -1046 2092 -1012 2268
rect 1012 2092 1046 2268
rect -1046 1656 -1012 1832
rect 1012 1656 1046 1832
rect -1046 1220 -1012 1396
rect 1012 1220 1046 1396
rect -1046 784 -1012 960
rect 1012 784 1046 960
rect -1046 348 -1012 524
rect 1012 348 1046 524
rect -1046 -88 -1012 88
rect 1012 -88 1046 88
rect -1046 -524 -1012 -348
rect 1012 -524 1046 -348
rect -1046 -960 -1012 -784
rect 1012 -960 1046 -784
rect -1046 -1396 -1012 -1220
rect 1012 -1396 1046 -1220
rect -1046 -1832 -1012 -1656
rect 1012 -1832 1046 -1656
rect -1046 -2268 -1012 -2092
rect 1012 -2268 1046 -2092
rect -1046 -2704 -1012 -2528
rect 1012 -2704 1046 -2528
rect -1046 -3140 -1012 -2964
rect 1012 -3140 1046 -2964
<< mvnsubdiff >>
rect -1192 3371 1192 3383
rect -1192 3337 -1084 3371
rect 1084 3337 1192 3371
rect -1192 3325 1192 3337
rect -1192 3275 -1134 3325
rect -1192 -3275 -1180 3275
rect -1146 -3275 -1134 3275
rect 1134 3275 1192 3325
rect -1192 -3325 -1134 -3275
rect 1134 -3275 1146 3275
rect 1180 -3275 1192 3275
rect 1134 -3325 1192 -3275
rect -1192 -3337 1192 -3325
rect -1192 -3371 -1084 -3337
rect 1084 -3371 1192 -3337
rect -1192 -3383 1192 -3371
<< mvnsubdiffcont >>
rect -1084 3337 1084 3371
rect -1180 -3275 -1146 3275
rect 1146 -3275 1180 3275
rect -1084 -3371 1084 -3337
<< poly >>
rect -1000 3233 1000 3249
rect -1000 3199 -984 3233
rect 984 3199 1000 3233
rect -1000 3152 1000 3199
rect -1000 2905 1000 2952
rect -1000 2871 -984 2905
rect 984 2871 1000 2905
rect -1000 2855 1000 2871
rect -1000 2797 1000 2813
rect -1000 2763 -984 2797
rect 984 2763 1000 2797
rect -1000 2716 1000 2763
rect -1000 2469 1000 2516
rect -1000 2435 -984 2469
rect 984 2435 1000 2469
rect -1000 2419 1000 2435
rect -1000 2361 1000 2377
rect -1000 2327 -984 2361
rect 984 2327 1000 2361
rect -1000 2280 1000 2327
rect -1000 2033 1000 2080
rect -1000 1999 -984 2033
rect 984 1999 1000 2033
rect -1000 1983 1000 1999
rect -1000 1925 1000 1941
rect -1000 1891 -984 1925
rect 984 1891 1000 1925
rect -1000 1844 1000 1891
rect -1000 1597 1000 1644
rect -1000 1563 -984 1597
rect 984 1563 1000 1597
rect -1000 1547 1000 1563
rect -1000 1489 1000 1505
rect -1000 1455 -984 1489
rect 984 1455 1000 1489
rect -1000 1408 1000 1455
rect -1000 1161 1000 1208
rect -1000 1127 -984 1161
rect 984 1127 1000 1161
rect -1000 1111 1000 1127
rect -1000 1053 1000 1069
rect -1000 1019 -984 1053
rect 984 1019 1000 1053
rect -1000 972 1000 1019
rect -1000 725 1000 772
rect -1000 691 -984 725
rect 984 691 1000 725
rect -1000 675 1000 691
rect -1000 617 1000 633
rect -1000 583 -984 617
rect 984 583 1000 617
rect -1000 536 1000 583
rect -1000 289 1000 336
rect -1000 255 -984 289
rect 984 255 1000 289
rect -1000 239 1000 255
rect -1000 181 1000 197
rect -1000 147 -984 181
rect 984 147 1000 181
rect -1000 100 1000 147
rect -1000 -147 1000 -100
rect -1000 -181 -984 -147
rect 984 -181 1000 -147
rect -1000 -197 1000 -181
rect -1000 -255 1000 -239
rect -1000 -289 -984 -255
rect 984 -289 1000 -255
rect -1000 -336 1000 -289
rect -1000 -583 1000 -536
rect -1000 -617 -984 -583
rect 984 -617 1000 -583
rect -1000 -633 1000 -617
rect -1000 -691 1000 -675
rect -1000 -725 -984 -691
rect 984 -725 1000 -691
rect -1000 -772 1000 -725
rect -1000 -1019 1000 -972
rect -1000 -1053 -984 -1019
rect 984 -1053 1000 -1019
rect -1000 -1069 1000 -1053
rect -1000 -1127 1000 -1111
rect -1000 -1161 -984 -1127
rect 984 -1161 1000 -1127
rect -1000 -1208 1000 -1161
rect -1000 -1455 1000 -1408
rect -1000 -1489 -984 -1455
rect 984 -1489 1000 -1455
rect -1000 -1505 1000 -1489
rect -1000 -1563 1000 -1547
rect -1000 -1597 -984 -1563
rect 984 -1597 1000 -1563
rect -1000 -1644 1000 -1597
rect -1000 -1891 1000 -1844
rect -1000 -1925 -984 -1891
rect 984 -1925 1000 -1891
rect -1000 -1941 1000 -1925
rect -1000 -1999 1000 -1983
rect -1000 -2033 -984 -1999
rect 984 -2033 1000 -1999
rect -1000 -2080 1000 -2033
rect -1000 -2327 1000 -2280
rect -1000 -2361 -984 -2327
rect 984 -2361 1000 -2327
rect -1000 -2377 1000 -2361
rect -1000 -2435 1000 -2419
rect -1000 -2469 -984 -2435
rect 984 -2469 1000 -2435
rect -1000 -2516 1000 -2469
rect -1000 -2763 1000 -2716
rect -1000 -2797 -984 -2763
rect 984 -2797 1000 -2763
rect -1000 -2813 1000 -2797
rect -1000 -2871 1000 -2855
rect -1000 -2905 -984 -2871
rect 984 -2905 1000 -2871
rect -1000 -2952 1000 -2905
rect -1000 -3199 1000 -3152
rect -1000 -3233 -984 -3199
rect 984 -3233 1000 -3199
rect -1000 -3249 1000 -3233
<< polycont >>
rect -984 3199 984 3233
rect -984 2871 984 2905
rect -984 2763 984 2797
rect -984 2435 984 2469
rect -984 2327 984 2361
rect -984 1999 984 2033
rect -984 1891 984 1925
rect -984 1563 984 1597
rect -984 1455 984 1489
rect -984 1127 984 1161
rect -984 1019 984 1053
rect -984 691 984 725
rect -984 583 984 617
rect -984 255 984 289
rect -984 147 984 181
rect -984 -181 984 -147
rect -984 -289 984 -255
rect -984 -617 984 -583
rect -984 -725 984 -691
rect -984 -1053 984 -1019
rect -984 -1161 984 -1127
rect -984 -1489 984 -1455
rect -984 -1597 984 -1563
rect -984 -1925 984 -1891
rect -984 -2033 984 -1999
rect -984 -2361 984 -2327
rect -984 -2469 984 -2435
rect -984 -2797 984 -2763
rect -984 -2905 984 -2871
rect -984 -3233 984 -3199
<< locali >>
rect -1180 3337 -1084 3371
rect 1084 3337 1180 3371
rect -1180 3275 -1146 3337
rect 1146 3275 1180 3337
rect -1000 3199 -984 3233
rect 984 3199 1000 3233
rect -1046 3140 -1012 3156
rect -1046 2948 -1012 2964
rect 1012 3140 1046 3156
rect 1012 2948 1046 2964
rect -1000 2871 -984 2905
rect 984 2871 1000 2905
rect -1000 2763 -984 2797
rect 984 2763 1000 2797
rect -1046 2704 -1012 2720
rect -1046 2512 -1012 2528
rect 1012 2704 1046 2720
rect 1012 2512 1046 2528
rect -1000 2435 -984 2469
rect 984 2435 1000 2469
rect -1000 2327 -984 2361
rect 984 2327 1000 2361
rect -1046 2268 -1012 2284
rect -1046 2076 -1012 2092
rect 1012 2268 1046 2284
rect 1012 2076 1046 2092
rect -1000 1999 -984 2033
rect 984 1999 1000 2033
rect -1000 1891 -984 1925
rect 984 1891 1000 1925
rect -1046 1832 -1012 1848
rect -1046 1640 -1012 1656
rect 1012 1832 1046 1848
rect 1012 1640 1046 1656
rect -1000 1563 -984 1597
rect 984 1563 1000 1597
rect -1000 1455 -984 1489
rect 984 1455 1000 1489
rect -1046 1396 -1012 1412
rect -1046 1204 -1012 1220
rect 1012 1396 1046 1412
rect 1012 1204 1046 1220
rect -1000 1127 -984 1161
rect 984 1127 1000 1161
rect -1000 1019 -984 1053
rect 984 1019 1000 1053
rect -1046 960 -1012 976
rect -1046 768 -1012 784
rect 1012 960 1046 976
rect 1012 768 1046 784
rect -1000 691 -984 725
rect 984 691 1000 725
rect -1000 583 -984 617
rect 984 583 1000 617
rect -1046 524 -1012 540
rect -1046 332 -1012 348
rect 1012 524 1046 540
rect 1012 332 1046 348
rect -1000 255 -984 289
rect 984 255 1000 289
rect -1000 147 -984 181
rect 984 147 1000 181
rect -1046 88 -1012 104
rect -1046 -104 -1012 -88
rect 1012 88 1046 104
rect 1012 -104 1046 -88
rect -1000 -181 -984 -147
rect 984 -181 1000 -147
rect -1000 -289 -984 -255
rect 984 -289 1000 -255
rect -1046 -348 -1012 -332
rect -1046 -540 -1012 -524
rect 1012 -348 1046 -332
rect 1012 -540 1046 -524
rect -1000 -617 -984 -583
rect 984 -617 1000 -583
rect -1000 -725 -984 -691
rect 984 -725 1000 -691
rect -1046 -784 -1012 -768
rect -1046 -976 -1012 -960
rect 1012 -784 1046 -768
rect 1012 -976 1046 -960
rect -1000 -1053 -984 -1019
rect 984 -1053 1000 -1019
rect -1000 -1161 -984 -1127
rect 984 -1161 1000 -1127
rect -1046 -1220 -1012 -1204
rect -1046 -1412 -1012 -1396
rect 1012 -1220 1046 -1204
rect 1012 -1412 1046 -1396
rect -1000 -1489 -984 -1455
rect 984 -1489 1000 -1455
rect -1000 -1597 -984 -1563
rect 984 -1597 1000 -1563
rect -1046 -1656 -1012 -1640
rect -1046 -1848 -1012 -1832
rect 1012 -1656 1046 -1640
rect 1012 -1848 1046 -1832
rect -1000 -1925 -984 -1891
rect 984 -1925 1000 -1891
rect -1000 -2033 -984 -1999
rect 984 -2033 1000 -1999
rect -1046 -2092 -1012 -2076
rect -1046 -2284 -1012 -2268
rect 1012 -2092 1046 -2076
rect 1012 -2284 1046 -2268
rect -1000 -2361 -984 -2327
rect 984 -2361 1000 -2327
rect -1000 -2469 -984 -2435
rect 984 -2469 1000 -2435
rect -1046 -2528 -1012 -2512
rect -1046 -2720 -1012 -2704
rect 1012 -2528 1046 -2512
rect 1012 -2720 1046 -2704
rect -1000 -2797 -984 -2763
rect 984 -2797 1000 -2763
rect -1000 -2905 -984 -2871
rect 984 -2905 1000 -2871
rect -1046 -2964 -1012 -2948
rect -1046 -3156 -1012 -3140
rect 1012 -2964 1046 -2948
rect 1012 -3156 1046 -3140
rect -1000 -3233 -984 -3199
rect 984 -3233 1000 -3199
rect -1180 -3337 -1146 -3275
rect 1146 -3337 1180 -3275
rect -1180 -3371 -1084 -3337
rect 1084 -3371 1180 -3337
<< viali >>
rect -984 3199 984 3233
rect -1046 2964 -1012 3140
rect 1012 2964 1046 3140
rect -984 2871 984 2905
rect -984 2763 984 2797
rect -1046 2528 -1012 2704
rect 1012 2528 1046 2704
rect -984 2435 984 2469
rect -984 2327 984 2361
rect -1046 2092 -1012 2268
rect 1012 2092 1046 2268
rect -984 1999 984 2033
rect -984 1891 984 1925
rect -1046 1656 -1012 1832
rect 1012 1656 1046 1832
rect -984 1563 984 1597
rect -984 1455 984 1489
rect -1046 1220 -1012 1396
rect 1012 1220 1046 1396
rect -984 1127 984 1161
rect -984 1019 984 1053
rect -1046 784 -1012 960
rect 1012 784 1046 960
rect -984 691 984 725
rect -984 583 984 617
rect -1046 348 -1012 524
rect 1012 348 1046 524
rect -984 255 984 289
rect -984 147 984 181
rect -1046 -88 -1012 88
rect 1012 -88 1046 88
rect -984 -181 984 -147
rect -984 -289 984 -255
rect -1046 -524 -1012 -348
rect 1012 -524 1046 -348
rect -984 -617 984 -583
rect -984 -725 984 -691
rect -1046 -960 -1012 -784
rect 1012 -960 1046 -784
rect -984 -1053 984 -1019
rect -984 -1161 984 -1127
rect -1046 -1396 -1012 -1220
rect 1012 -1396 1046 -1220
rect -984 -1489 984 -1455
rect -984 -1597 984 -1563
rect -1046 -1832 -1012 -1656
rect 1012 -1832 1046 -1656
rect -984 -1925 984 -1891
rect -984 -2033 984 -1999
rect -1046 -2268 -1012 -2092
rect 1012 -2268 1046 -2092
rect -984 -2361 984 -2327
rect -984 -2469 984 -2435
rect -1046 -2704 -1012 -2528
rect 1012 -2704 1046 -2528
rect -984 -2797 984 -2763
rect -984 -2905 984 -2871
rect -1046 -3140 -1012 -2964
rect 1012 -3140 1046 -2964
rect -984 -3233 984 -3199
<< metal1 >>
rect -996 3233 996 3239
rect -996 3199 -984 3233
rect 984 3199 996 3233
rect -996 3193 996 3199
rect -1052 3140 -1006 3152
rect -1052 2964 -1046 3140
rect -1012 2964 -1006 3140
rect -1052 2952 -1006 2964
rect 1006 3140 1052 3152
rect 1006 2964 1012 3140
rect 1046 2964 1052 3140
rect 1006 2952 1052 2964
rect -996 2905 996 2911
rect -996 2871 -984 2905
rect 984 2871 996 2905
rect -996 2865 996 2871
rect -996 2797 996 2803
rect -996 2763 -984 2797
rect 984 2763 996 2797
rect -996 2757 996 2763
rect -1052 2704 -1006 2716
rect -1052 2528 -1046 2704
rect -1012 2528 -1006 2704
rect -1052 2516 -1006 2528
rect 1006 2704 1052 2716
rect 1006 2528 1012 2704
rect 1046 2528 1052 2704
rect 1006 2516 1052 2528
rect -996 2469 996 2475
rect -996 2435 -984 2469
rect 984 2435 996 2469
rect -996 2429 996 2435
rect -996 2361 996 2367
rect -996 2327 -984 2361
rect 984 2327 996 2361
rect -996 2321 996 2327
rect -1052 2268 -1006 2280
rect -1052 2092 -1046 2268
rect -1012 2092 -1006 2268
rect -1052 2080 -1006 2092
rect 1006 2268 1052 2280
rect 1006 2092 1012 2268
rect 1046 2092 1052 2268
rect 1006 2080 1052 2092
rect -996 2033 996 2039
rect -996 1999 -984 2033
rect 984 1999 996 2033
rect -996 1993 996 1999
rect -996 1925 996 1931
rect -996 1891 -984 1925
rect 984 1891 996 1925
rect -996 1885 996 1891
rect -1052 1832 -1006 1844
rect -1052 1656 -1046 1832
rect -1012 1656 -1006 1832
rect -1052 1644 -1006 1656
rect 1006 1832 1052 1844
rect 1006 1656 1012 1832
rect 1046 1656 1052 1832
rect 1006 1644 1052 1656
rect -996 1597 996 1603
rect -996 1563 -984 1597
rect 984 1563 996 1597
rect -996 1557 996 1563
rect -996 1489 996 1495
rect -996 1455 -984 1489
rect 984 1455 996 1489
rect -996 1449 996 1455
rect -1052 1396 -1006 1408
rect -1052 1220 -1046 1396
rect -1012 1220 -1006 1396
rect -1052 1208 -1006 1220
rect 1006 1396 1052 1408
rect 1006 1220 1012 1396
rect 1046 1220 1052 1396
rect 1006 1208 1052 1220
rect -996 1161 996 1167
rect -996 1127 -984 1161
rect 984 1127 996 1161
rect -996 1121 996 1127
rect -996 1053 996 1059
rect -996 1019 -984 1053
rect 984 1019 996 1053
rect -996 1013 996 1019
rect -1052 960 -1006 972
rect -1052 784 -1046 960
rect -1012 784 -1006 960
rect -1052 772 -1006 784
rect 1006 960 1052 972
rect 1006 784 1012 960
rect 1046 784 1052 960
rect 1006 772 1052 784
rect -996 725 996 731
rect -996 691 -984 725
rect 984 691 996 725
rect -996 685 996 691
rect -996 617 996 623
rect -996 583 -984 617
rect 984 583 996 617
rect -996 577 996 583
rect -1052 524 -1006 536
rect -1052 348 -1046 524
rect -1012 348 -1006 524
rect -1052 336 -1006 348
rect 1006 524 1052 536
rect 1006 348 1012 524
rect 1046 348 1052 524
rect 1006 336 1052 348
rect -996 289 996 295
rect -996 255 -984 289
rect 984 255 996 289
rect -996 249 996 255
rect -996 181 996 187
rect -996 147 -984 181
rect 984 147 996 181
rect -996 141 996 147
rect -1052 88 -1006 100
rect -1052 -88 -1046 88
rect -1012 -88 -1006 88
rect -1052 -100 -1006 -88
rect 1006 88 1052 100
rect 1006 -88 1012 88
rect 1046 -88 1052 88
rect 1006 -100 1052 -88
rect -996 -147 996 -141
rect -996 -181 -984 -147
rect 984 -181 996 -147
rect -996 -187 996 -181
rect -996 -255 996 -249
rect -996 -289 -984 -255
rect 984 -289 996 -255
rect -996 -295 996 -289
rect -1052 -348 -1006 -336
rect -1052 -524 -1046 -348
rect -1012 -524 -1006 -348
rect -1052 -536 -1006 -524
rect 1006 -348 1052 -336
rect 1006 -524 1012 -348
rect 1046 -524 1052 -348
rect 1006 -536 1052 -524
rect -996 -583 996 -577
rect -996 -617 -984 -583
rect 984 -617 996 -583
rect -996 -623 996 -617
rect -996 -691 996 -685
rect -996 -725 -984 -691
rect 984 -725 996 -691
rect -996 -731 996 -725
rect -1052 -784 -1006 -772
rect -1052 -960 -1046 -784
rect -1012 -960 -1006 -784
rect -1052 -972 -1006 -960
rect 1006 -784 1052 -772
rect 1006 -960 1012 -784
rect 1046 -960 1052 -784
rect 1006 -972 1052 -960
rect -996 -1019 996 -1013
rect -996 -1053 -984 -1019
rect 984 -1053 996 -1019
rect -996 -1059 996 -1053
rect -996 -1127 996 -1121
rect -996 -1161 -984 -1127
rect 984 -1161 996 -1127
rect -996 -1167 996 -1161
rect -1052 -1220 -1006 -1208
rect -1052 -1396 -1046 -1220
rect -1012 -1396 -1006 -1220
rect -1052 -1408 -1006 -1396
rect 1006 -1220 1052 -1208
rect 1006 -1396 1012 -1220
rect 1046 -1396 1052 -1220
rect 1006 -1408 1052 -1396
rect -996 -1455 996 -1449
rect -996 -1489 -984 -1455
rect 984 -1489 996 -1455
rect -996 -1495 996 -1489
rect -996 -1563 996 -1557
rect -996 -1597 -984 -1563
rect 984 -1597 996 -1563
rect -996 -1603 996 -1597
rect -1052 -1656 -1006 -1644
rect -1052 -1832 -1046 -1656
rect -1012 -1832 -1006 -1656
rect -1052 -1844 -1006 -1832
rect 1006 -1656 1052 -1644
rect 1006 -1832 1012 -1656
rect 1046 -1832 1052 -1656
rect 1006 -1844 1052 -1832
rect -996 -1891 996 -1885
rect -996 -1925 -984 -1891
rect 984 -1925 996 -1891
rect -996 -1931 996 -1925
rect -996 -1999 996 -1993
rect -996 -2033 -984 -1999
rect 984 -2033 996 -1999
rect -996 -2039 996 -2033
rect -1052 -2092 -1006 -2080
rect -1052 -2268 -1046 -2092
rect -1012 -2268 -1006 -2092
rect -1052 -2280 -1006 -2268
rect 1006 -2092 1052 -2080
rect 1006 -2268 1012 -2092
rect 1046 -2268 1052 -2092
rect 1006 -2280 1052 -2268
rect -996 -2327 996 -2321
rect -996 -2361 -984 -2327
rect 984 -2361 996 -2327
rect -996 -2367 996 -2361
rect -996 -2435 996 -2429
rect -996 -2469 -984 -2435
rect 984 -2469 996 -2435
rect -996 -2475 996 -2469
rect -1052 -2528 -1006 -2516
rect -1052 -2704 -1046 -2528
rect -1012 -2704 -1006 -2528
rect -1052 -2716 -1006 -2704
rect 1006 -2528 1052 -2516
rect 1006 -2704 1012 -2528
rect 1046 -2704 1052 -2528
rect 1006 -2716 1052 -2704
rect -996 -2763 996 -2757
rect -996 -2797 -984 -2763
rect 984 -2797 996 -2763
rect -996 -2803 996 -2797
rect -996 -2871 996 -2865
rect -996 -2905 -984 -2871
rect 984 -2905 996 -2871
rect -996 -2911 996 -2905
rect -1052 -2964 -1006 -2952
rect -1052 -3140 -1046 -2964
rect -1012 -3140 -1006 -2964
rect -1052 -3152 -1006 -3140
rect 1006 -2964 1052 -2952
rect 1006 -3140 1012 -2964
rect 1046 -3140 1052 -2964
rect 1006 -3152 1052 -3140
rect -996 -3199 996 -3193
rect -996 -3233 -984 -3199
rect 984 -3233 996 -3199
rect -996 -3239 996 -3233
<< properties >>
string FIXED_BBOX -1163 -3354 1163 3354
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
