magic
tech sky130A
timestamp 1717294357
<< metal1 >>
rect 4582 -2684 4609 -2681
rect 4582 -2888 4609 -2884
<< via1 >>
rect 4582 -2884 4609 -2684
<< metal2 >>
rect 4579 -2884 4582 -2684
rect 4609 -2884 4612 -2684
<< end >>
