magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< pwell >>
rect -2228 -363 2228 363
<< mvnmos >>
rect -2000 -105 2000 105
<< mvndiff >>
rect -2058 93 -2000 105
rect -2058 -93 -2046 93
rect -2012 -93 -2000 93
rect -2058 -105 -2000 -93
rect 2000 93 2058 105
rect 2000 -93 2012 93
rect 2046 -93 2058 93
rect 2000 -105 2058 -93
<< mvndiffc >>
rect -2046 -93 -2012 93
rect 2012 -93 2046 93
<< mvpsubdiff >>
rect -2192 315 2192 327
rect -2192 281 -2084 315
rect 2084 281 2192 315
rect -2192 269 2192 281
rect -2192 219 -2134 269
rect -2192 -219 -2180 219
rect -2146 -219 -2134 219
rect 2134 219 2192 269
rect -2192 -269 -2134 -219
rect 2134 -219 2146 219
rect 2180 -219 2192 219
rect 2134 -269 2192 -219
rect -2192 -281 2192 -269
rect -2192 -315 -2084 -281
rect 2084 -315 2192 -281
rect -2192 -327 2192 -315
<< mvpsubdiffcont >>
rect -2084 281 2084 315
rect -2180 -219 -2146 219
rect 2146 -219 2180 219
rect -2084 -315 2084 -281
<< poly >>
rect -2000 177 2000 193
rect -2000 143 -1984 177
rect 1984 143 2000 177
rect -2000 105 2000 143
rect -2000 -143 2000 -105
rect -2000 -177 -1984 -143
rect 1984 -177 2000 -143
rect -2000 -193 2000 -177
<< polycont >>
rect -1984 143 1984 177
rect -1984 -177 1984 -143
<< locali >>
rect -2180 281 -2084 315
rect 2084 281 2180 315
rect -2180 219 -2146 281
rect 2146 219 2180 281
rect -2000 143 -1984 177
rect 1984 143 2000 177
rect -2046 93 -2012 109
rect -2046 -109 -2012 -93
rect 2012 93 2046 109
rect 2012 -109 2046 -93
rect -2000 -177 -1984 -143
rect 1984 -177 2000 -143
rect -2180 -281 -2146 -219
rect 2146 -281 2180 -219
rect -2180 -315 -2084 -281
rect 2084 -315 2180 -281
<< viali >>
rect -1984 143 1984 177
rect -2046 -93 -2012 93
rect 2012 -93 2046 93
rect -1984 -177 1984 -143
<< metal1 >>
rect -1996 177 1996 183
rect -1996 143 -1984 177
rect 1984 143 1996 177
rect -1996 137 1996 143
rect -2052 93 -2006 105
rect -2052 -93 -2046 93
rect -2012 -93 -2006 93
rect -2052 -105 -2006 -93
rect 2006 93 2052 105
rect 2006 -93 2012 93
rect 2046 -93 2052 93
rect 2006 -105 2052 -93
rect -1996 -143 1996 -137
rect -1996 -177 -1984 -143
rect 1984 -177 1996 -143
rect -1996 -183 1996 -177
<< properties >>
string FIXED_BBOX -2163 -298 2163 298
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.05 l 20.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
