magic
tech sky130A
timestamp 1717294357
<< metal1 >>
rect 8313 -3180 8382 -3177
rect 8313 -3243 8316 -3180
rect 8379 -3243 8382 -3180
rect 8313 -3246 8382 -3243
<< via1 >>
rect 8316 -3243 8379 -3180
<< metal2 >>
rect 8313 -3180 8382 -3177
rect 8313 -3243 8316 -3180
rect 8379 -3243 8382 -3180
rect 8313 -3246 8382 -3243
<< end >>
