* NGSPICE file created from sky130_am_ip__ldo_01v8.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BWAZV5 a_n700_n197# a_700_n100# w_n958_n397#
+ a_n758_n100#
X0 a_700_n100# a_n700_n197# a_n758_n100# w_n958_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_A2FZRM a_n900_n188# a_n900_n1024# a_900_n518#
+ a_n900_648# a_n958_318# a_n958_n518# a_900_736# a_n1102_n1158# a_900_n100# a_900_n936#
+ a_900_318# a_n900_230# a_n958_n100# a_n958_736# a_n958_n936# a_n900_n606#
X0 a_900_n100# a_n900_n188# a_n958_n100# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X1 a_900_n518# a_n900_n606# a_n958_n518# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X2 a_900_318# a_n900_230# a_n958_318# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X3 a_900_n936# a_n900_n1024# a_n958_n936# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X4 a_900_736# a_n900_648# a_n958_736# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6 a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PC2PN5 w_n1258_n397# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1258_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.12188 ps=1.075 w=0.75 l=0.5
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X12 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.12188 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69K6TN a_700_n100# a_n758_n100# a_n700_n188#
+ a_n902_n322#
X0 a_700_n100# a_n700_n188# a_n758_n100# a_n902_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QZEXQH a_1044_n1416# a_214_n1416# a_n1114_n1416#
+ a_546_984# a_n1114_984# a_n118_984# a_48_n1416# a_1376_n1416# a_n450_984# a_n782_n1416#
+ a_878_984# a_546_n1416# a_n1446_984# a_712_984# a_n1446_n1416# a_n284_n1416# a_n616_n1416#
+ a_n782_984# a_1210_n1416# a_1044_984# a_878_n1416# a_n118_n1416# a_n616_984# a_48_984#
+ a_380_984# a_1376_984# a_n948_n1416# a_n1576_n1546# a_380_n1416# a_n948_984# a_712_n1416#
+ a_1210_984# a_214_984# a_n1280_n1416# a_n284_984# a_n450_n1416# a_n1280_984#
X0 a_n118_984# a_n118_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n1280_984# a_n1280_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_n948_984# a_n948_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_1210_984# a_1210_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n616_984# a_n616_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_380_984# a_380_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_878_984# a_878_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_546_984# a_546_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n1446_984# a_n1446_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_214_984# a_214_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_1376_984# a_1376_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n1114_984# a_n1114_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_n284_984# a_n284_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_1044_984# a_1044_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_n450_984# a_n450_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_48_984# a_48_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_712_984# a_712_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_n782_984# a_n782_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H a_1044_n1416# a_214_n1416# a_n2276_984#
+ a_n2110_n1416# a_1542_984# a_n1114_n1416# a_2870_n1416# a_546_984# a_n1114_984#
+ a_n118_984# a_n2110_984# a_1874_n1416# a_2538_984# a_48_n1416# a_n2940_n1416# a_2372_n1416#
+ a_n1944_n1416# a_1874_984# a_n782_n1416# a_n450_984# a_1376_n1416# a_2870_984# a_878_984#
+ a_2704_n1416# a_546_n1416# a_n1446_984# a_n2442_984# a_1708_n1416# a_n2442_n1416#
+ a_n1446_n1416# a_712_984# a_n284_n1416# a_1708_984# a_2206_n1416# a_2704_984# a_n782_984#
+ a_n616_n1416# a_n1778_984# a_n2774_984# a_1210_n1416# a_1044_984# a_2040_984# a_n1612_984#
+ a_878_n1416# a_n118_n1416# a_n616_984# a_n2774_n1416# a_n2608_984# a_n1778_n1416#
+ a_48_984# a_2538_n1416# a_380_984# a_1376_984# a_n948_n1416# a_2372_984# a_n1944_984#
+ a_380_n1416# a_n2276_n1416# a_n948_984# a_n3070_n1546# a_n2940_984# a_1542_n1416#
+ a_712_n1416# a_n2608_n1416# a_1210_984# a_n1280_n1416# a_214_984# a_2040_n1416#
+ a_n1612_n1416# a_n1280_984# a_2206_984# a_n450_n1416# a_n284_984#
X0 a_n2276_984# a_n2276_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n118_984# a_n118_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_1542_984# a_1542_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n1280_984# a_n1280_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n948_984# a_n948_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_2704_984# a_2704_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_1210_984# a_1210_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_1708_984# a_1708_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n616_984# a_n616_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_380_984# a_380_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_n2774_984# a_n2774_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n2110_984# a_n2110_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_878_984# a_878_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_n1778_984# a_n1778_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_n2442_984# a_n2442_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_n2940_984# a_n2940_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_546_984# a_546_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_n1446_984# a_n1446_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X18 a_2372_984# a_2372_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X19 a_214_984# a_214_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X20 a_1376_984# a_1376_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X21 a_n2608_984# a_n2608_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X22 a_n1114_984# a_n1114_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X23 a_n284_984# a_n284_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X24 a_2040_984# a_2040_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X25 a_2538_984# a_2538_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X26 a_1044_984# a_1044_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X27 a_n1944_984# a_n1944_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X28 a_n450_984# a_n450_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X29 a_48_984# a_48_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X30 a_2206_984# a_2206_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X31 a_2870_984# a_2870_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X32 a_712_984# a_712_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X33 a_1874_984# a_1874_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X34 a_n1612_984# a_n1612_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X35 a_n782_984# a_n782_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_743D3R a_n248_n2546# a_48_n2416# a_n118_1984#
+ a_n118_n2416# a_48_1984#
X0 a_48_1984# a_48_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X1 a_n118_1984# a_n118_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MRZGNS c1_n1646_n1500# m3_n1686_n1540#
X0 c1_n1646_n1500# m3_n1686_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PXBJUB a_n1000_n188# a_n1192_n322# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1192_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_47NWVV a_n258_n100# a_n200_n197# a_200_n100#
+ w_n458_n397#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n458_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YHRXVR a_n129_n2415# a_819_2457# a_n977_2545#
+ a_n1609_n4763# a_n1135_n1109# a_n1551_21# a_n503_n4763# a_603_n3545# a_1235_109#
+ a_n1609_n1109# a_n29_4981# a_445_3763# a_n1135_109# a_n1077_2457# a_n1235_n2415#
+ a_n503_n1109# a_1393_4981# a_n29_1327# a_345_2457# a_1235_n3545# a_977_n3633# a_n761_3675#
+ a_n603_n2415# a_1393_1327# a_1293_3675# a_n919_2457# a_977_21# a_n345_n4763# a_445_n3545#
+ a_n503_2545# a_129_2545# a_n1077_n2415# a_n187_4981# a_n1293_2545# a_n819_n4763#
+ a_919_n3545# a_n345_n1109# a_n1551_3675# a_187_21# a_1077_3763# a_n1451_n4763# a_29_n4851#
+ a_1077_n3545# a_977_2457# a_n187_1327# a_n819_n1109# a_503_n2415# a_n129_n1197#
+ a_n445_n2415# a_n445_2457# a_n1451_n1109# a_n977_109# a_1077_109# a_n919_n2415#
+ a_n1235_n1197# a_1135_n2415# a_n1551_n2415# a_29_4893# a_n187_n4763# a_287_n3545#
+ a_1451_21# a_29_1239# a_1551_n3545# a_n187_n1109# a_603_3763# a_n603_n1197# a_n1293_n4763#
+ a_n1235_2457# a_n129_4893# a_345_n2415# a_1551_4981# a_n287_n2415# a_129_109# a_n1293_n1109#
+ a_n129_1239# a_503_2457# a_n661_2545# a_n445_21# a_819_n2415# a_29_n6069# a_287_2545#
+ a_n661_n4763# a_761_n3545# a_1551_1327# a_n819_4981# a_n29_n3545# a_187_4893# a_1451_3675#
+ a_n1077_n1197# a_n1393_n2415# a_n661_n1109# a_n819_1327# a_187_1239# a_1393_n3545#
+ a_503_n1197# a_n445_n1197# a_n761_n2415# a_n345_4981# a_n1451_2545# a_187_n2415#
+ a_n919_n1197# a_n1609_109# a_n1609_4981# a_1235_3763# a_1135_n1197# a_n345_1327#
+ a_n1551_n1197# a_1451_n2415# a_n603_2457# a_n1609_1327# a_129_n5981# a_1135_2457#
+ a_n1077_21# a_761_3763# a_n977_n4763# a_n1393_2457# a_n287_4893# a_129_n2327# a_345_n1197#
+ a_n1135_4981# a_n977_n1109# a_661_n2415# a_n287_1239# a_661_2457# a_n29_109# a_n287_n1197#
+ a_919_2545# a_1551_109# a_819_n1197# a_n129_n4851# a_819_4893# a_n1135_1327# a_n977_4981#
+ a_n1451_109# a_n1135_n3545# a_345_21# a_29_21# a_n1393_n1197# a_1293_n2415# a_603_n5981#
+ a_819_1239# a_n977_1327# a_n1609_n3545# a_n1077_4893# a_n1235_n4851# a_603_n2327#
+ a_n503_n3545# a_n29_3763# a_445_2545# a_n1077_1239# a_n503_109# a_n761_n1197# a_1235_n5981#
+ a_345_4893# a_187_n1197# a_1393_3763# a_n603_n4851# a_603_109# a_345_1239# a_1235_n2327#
+ a_1451_n1197# a_977_n2415# a_n761_2457# a_1293_2457# a_n919_4893# a_n503_4981# a_445_n5981#
+ a_129_4981# a_n1077_n4851# a_n129_n6069# a_n1293_4981# a_n919_1239# a_919_n5981#
+ a_n503_1327# a_n603_21# a_445_n2327# a_n345_n3545# a_661_n1197# a_129_1327# a_1077_n5981#
+ a_n187_3763# a_n1293_1327# a_1393_109# a_n819_n3545# a_977_4893# a_919_n2327# a_503_n4851#
+ a_n1293_109# a_n1235_n6069# a_n445_n4851# a_n1551_2457# a_1077_2545# a_n445_4893#
+ a_29_n3633# a_n1451_n3545# a_1077_n2327# a_977_1239# a_1293_n1197# a_n919_n4851#
+ a_n445_1239# a_1135_n4851# a_n1551_n4851# a_n603_n6069# a_287_n5981# a_n345_109#
+ a_29_3675# a_1551_n5981# a_287_n2327# a_n187_n3545# a_445_109# a_n1235_4893# a_1551_n2327#
+ a_345_n4851# a_977_n1197# a_n1077_n6069# a_n287_n4851# a_n1235_21# a_603_2545# a_n129_3675#
+ a_n1235_1239# a_n1293_n3545# a_503_4893# a_n661_4981# a_819_n4851# a_287_4981# a_761_n5981#
+ a_1551_3763# a_n29_n5981# a_503_n6069# a_503_1239# a_n661_1327# a_n1393_n4851# a_n445_n6069#
+ a_287_1327# a_761_n2327# a_n661_n3545# a_n819_3763# a_187_3675# a_n29_n2327# a_1451_2457#
+ a_503_21# a_n919_n6069# a_1393_n5981# a_1135_n6069# a_n1551_n6069# a_n761_n4851#
+ a_n1451_4981# a_1393_n2327# a_187_n4851# a_n345_3763# a_n1451_1327# a_1451_n4851#
+ a_n187_109# a_n1609_3763# a_1235_2545# a_n603_4893# a_345_n6069# a_n287_n6069# a_1135_4893#
+ a_287_109# a_n1393_4893# a_819_n6069# a_n603_1239# a_129_n4763# a_1135_1239# a_761_2545#
+ a_n977_n3545# a_661_n4851# a_n287_3675# a_n1393_1239# a_n1393_n6069# a_661_4893#
+ a_919_4981# a_129_n1109# a_n1135_3763# a_n1135_n5981# a_661_1239# a_919_1327# a_n129_n3633#
+ a_1293_n4851# a_819_3675# a_n977_3763# a_n1609_n5981# a_n761_n6069# a_n1135_n2327#
+ a_1135_21# a_187_n6069# a_n503_n5981# a_603_n4763# a_n919_21# a_n1609_n2327# a_445_4981#
+ a_n1077_3675# a_n1235_n3633# a_1451_n6069# a_603_n1109# a_n503_n2327# a_n761_21#
+ a_n1753_n6203# a_n29_2545# a_445_1327# a_345_3675# a_n129_21# a_1235_n4763# a_977_n4851#
+ a_n603_n3633# a_n761_4893# a_1393_2545# a_n819_109# a_1293_4893# a_1235_n1109# a_661_n6069#
+ a_919_109# a_n761_1239# a_1293_1239# a_n919_3675# a_n345_n5981# a_n503_3763# a_445_n4763#
+ a_129_3763# a_n1077_n3633# a_1293_n6069# a_n1293_3763# a_n819_n5981# a_919_n4763#
+ a_445_n1109# a_n345_n2327# a_1077_4981# a_n1551_4893# a_n1451_n5981# a_1077_n4763#
+ a_977_3675# a_n187_2545# a_919_n1109# a_n819_n2327# a_503_n3633# a_n445_n3633# a_n661_109#
+ a_n445_3675# a_n1551_1239# a_1077_1327# a_n1393_21# a_29_n2415# a_n1451_n2327# a_1077_n1109#
+ a_761_109# a_n919_n3633# a_1135_n3633# a_n1551_n3633# a_977_n6069# a_819_21# a_n187_n5981#
+ a_287_n4763# a_661_21# a_29_2457# a_n187_n2327# a_1551_n4763# a_287_n1109# a_603_4981#
+ a_n1235_3675# a_n1293_n5981# a_345_n3633# a_1551_n1109# a_n287_n3633# a_603_1327#
+ a_n129_2457# a_n1293_n2327# a_503_3675# a_n661_3763# a_819_n3633# a_287_3763# a_n661_n5981#
+ a_761_n4763# a_1551_2545# a_n29_n4763# a_1451_4893# a_n1393_n3633# a_n661_n2327#
+ a_761_n1109# a_n819_2545# a_187_2457# a_1451_1239# a_n29_n1109# a_1393_n4763# a_n761_n3633#
+ a_29_n1197# a_n1451_3763# a_187_n3633# a_1393_n1109# a_1235_4981# a_1451_n3633#
+ a_n345_2545# a_n603_3675# a_n1609_2545# a_1235_1327# a_1293_21# a_1135_3675# a_761_4981#
+ a_n977_n5981# a_n1393_3675# a_129_n3545# a_761_1327# a_n977_n2327# a_661_n3633#
+ a_n287_2457# a_661_3675# a_919_3763# a_n287_21# a_n1135_2545# a_n1135_n4763# a_1293_n3633#
X0 a_n661_109# a_n761_21# a_n819_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_n187_n4763# a_n287_n4851# a_n345_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X2 a_1551_n5981# a_1451_n6069# a_1393_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X3 a_n29_n5981# a_n129_n6069# a_n187_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X4 a_129_n2327# a_29_n2415# a_n29_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X5 a_761_4981# a_661_4893# a_603_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X6 a_1393_2545# a_1293_2457# a_1235_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X7 a_n187_4981# a_n287_4893# a_n345_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X8 a_n1293_2545# a_n1393_2457# a_n1451_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X9 a_129_109# a_29_21# a_n29_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X10 a_445_n1109# a_345_n1197# a_287_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X11 a_287_3763# a_187_3675# a_129_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X12 a_n187_109# a_n287_21# a_n345_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X13 a_n187_n5981# a_n287_n6069# a_n345_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X14 a_129_n3545# a_29_n3633# a_n29_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X15 a_n1293_3763# a_n1393_3675# a_n1451_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X16 a_1393_3763# a_1293_3675# a_1235_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X17 a_n345_1327# a_n445_1239# a_n503_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X18 a_445_n2327# a_345_n2415# a_287_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X19 a_287_4981# a_187_4893# a_129_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X20 a_919_n1109# a_819_n1197# a_761_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X21 a_n819_109# a_n919_21# a_n977_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X22 a_129_n4763# a_29_n4851# a_n29_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X23 a_n1293_4981# a_n1393_4893# a_n1451_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X24 a_1393_4981# a_1293_4893# a_1235_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X25 a_129_1327# a_29_1239# a_n29_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X26 a_n345_109# a_n445_21# a_n503_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X27 a_n345_2545# a_n445_2457# a_n503_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X28 a_445_n3545# a_345_n3633# a_287_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X29 a_445_1327# a_345_1239# a_287_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X30 a_n1451_n1109# a_n1551_n1197# a_n1609_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X31 a_919_n2327# a_819_n2415# a_761_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X32 a_1077_n1109# a_977_n1197# a_919_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X33 a_129_n5981# a_29_n6069# a_n29_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X34 a_129_2545# a_29_2457# a_n29_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X35 a_n345_3763# a_n445_3675# a_n503_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X36 a_n1451_1327# a_n1551_1239# a_n1609_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X37 a_1551_1327# a_1451_1239# a_1393_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X38 a_445_n4763# a_345_n4851# a_287_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X39 a_n503_109# a_n603_21# a_n661_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X40 a_445_2545# a_345_2457# a_287_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X41 a_919_n3545# a_819_n3633# a_761_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X42 a_1077_n2327# a_977_n2415# a_919_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X43 a_n1451_n2327# a_n1551_n2415# a_n1609_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X44 a_n345_n1109# a_n445_n1197# a_n503_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X45 a_129_3763# a_29_3675# a_n29_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X46 a_1551_2545# a_1451_2457# a_1393_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X47 a_n345_4981# a_n445_4893# a_n503_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X48 a_n1451_2545# a_n1551_2457# a_n1609_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X49 a_445_n5981# a_345_n6069# a_287_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X50 a_n29_109# a_n129_21# a_n187_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X51 a_445_3763# a_345_3675# a_287_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X52 a_n977_1327# a_n1077_1239# a_n1135_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X53 a_919_n4763# a_819_n4851# a_761_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X54 a_1077_n3545# a_977_n3633# a_919_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X55 a_n1451_n3545# a_n1551_n3633# a_n1609_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X56 a_n345_n2327# a_n445_n2415# a_n503_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X57 a_129_4981# a_29_4893# a_n29_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X58 a_1551_3763# a_1451_3675# a_1393_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X59 a_1077_1327# a_977_1239# a_919_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X60 a_n1451_3763# a_n1551_3675# a_n1609_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X61 a_1393_109# a_1293_21# a_1235_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X62 a_n503_1327# a_n603_1239# a_n661_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X63 a_n819_n1109# a_n919_n1197# a_n977_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X64 a_445_4981# a_345_4893# a_287_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X65 a_n977_2545# a_n1077_2457# a_n1135_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X66 a_919_n5981# a_819_n6069# a_761_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X67 a_1077_n4763# a_977_n4851# a_919_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X68 a_n1451_n4763# a_n1551_n4851# a_n1609_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X69 a_1077_109# a_977_21# a_919_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X70 a_n977_n1109# a_n1077_n1197# a_n1135_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X71 a_n345_n3545# a_n445_n3633# a_n503_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X72 a_1551_4981# a_1451_4893# a_1393_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X73 a_1077_2545# a_977_2457# a_919_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X74 a_n1451_4981# a_n1551_4893# a_n1609_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X75 a_1235_n1109# a_1135_n1197# a_1077_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X76 a_n503_2545# a_n603_2457# a_n661_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X77 a_1551_109# a_1451_21# a_1393_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X78 a_n819_n2327# a_n919_n2415# a_n977_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X79 a_n977_3763# a_n1077_3675# a_n1135_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X80 a_1077_n5981# a_977_n6069# a_919_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X81 a_n1451_n5981# a_n1551_n6069# a_n1609_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X82 a_n29_1327# a_n129_1239# a_n187_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X83 a_603_1327# a_503_1239# a_445_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X84 a_n977_n2327# a_n1077_n2415# a_n1135_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X85 a_n345_n4763# a_n445_n4851# a_n503_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X86 a_1077_3763# a_977_3675# a_919_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X87 a_1235_n2327# a_1135_n2415# a_1077_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X88 a_1393_n1109# a_1293_n1197# a_1235_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X89 a_n503_3763# a_n603_3675# a_n661_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X90 a_761_109# a_661_21# a_603_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X91 a_n819_n3545# a_n919_n3633# a_n977_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X92 a_603_n1109# a_503_n1197# a_445_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X93 a_n977_4981# a_n1077_4893# a_n1135_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X94 a_n29_2545# a_n129_2457# a_n187_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X95 a_603_2545# a_503_2457# a_445_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X96 a_n977_n3545# a_n1077_n3633# a_n1135_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X97 a_n345_n5981# a_n445_n6069# a_n503_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X98 a_1077_4981# a_977_4893# a_919_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X99 a_1235_n3545# a_1135_n3633# a_1077_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X100 a_1393_n2327# a_1293_n2415# a_1235_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X101 a_n503_4981# a_n603_4893# a_n661_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X102 a_287_109# a_187_21# a_129_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X103 a_n819_n4763# a_n919_n4851# a_n977_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X104 a_603_n2327# a_503_n2415# a_445_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X105 a_761_n1109# a_661_n1197# a_603_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X106 a_1235_1327# a_1135_1239# a_1077_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X107 a_1235_109# a_1135_21# a_1077_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X108 a_n29_3763# a_n129_3675# a_n187_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X109 a_603_3763# a_503_3675# a_445_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X110 a_n1135_1327# a_n1235_1239# a_n1293_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X111 a_n977_n4763# a_n1077_n4851# a_n1135_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X112 a_1235_n4763# a_1135_n4851# a_1077_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X113 a_1393_n3545# a_1293_n3633# a_1235_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X114 a_919_109# a_819_21# a_761_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X115 a_n819_n5981# a_n919_n6069# a_n977_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X116 a_603_n3545# a_503_n3633# a_445_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X117 a_761_n2327# a_661_n2415# a_603_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X118 a_1235_2545# a_1135_2457# a_1077_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X119 a_445_109# a_345_21# a_287_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X120 a_n29_4981# a_n129_4893# a_n187_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X121 a_603_4981# a_503_4893# a_445_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X122 a_n1135_2545# a_n1235_2457# a_n1293_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X123 a_n977_n5981# a_n1077_n6069# a_n1135_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X124 a_1235_n5981# a_1135_n6069# a_1077_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X125 a_1393_n4763# a_1293_n4851# a_1235_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X126 a_761_n3545# a_661_n3633# a_603_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X127 a_603_n4763# a_503_n4851# a_445_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X128 a_1235_3763# a_1135_3675# a_1077_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X129 a_n1135_3763# a_n1235_3675# a_n1293_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X130 a_603_109# a_503_21# a_445_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X131 a_1393_n5981# a_1293_n6069# a_1235_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X132 a_n503_n1109# a_n603_n1197# a_n661_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X133 a_761_n4763# a_661_n4851# a_603_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X134 a_603_n5981# a_503_n6069# a_445_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X135 a_287_n1109# a_187_n1197# a_129_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X136 a_1235_4981# a_1135_4893# a_1077_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X137 a_n1135_4981# a_n1235_4893# a_n1293_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X138 a_n661_n1109# a_n761_n1197# a_n819_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X139 a_n503_n2327# a_n603_n2415# a_n661_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X140 a_761_n5981# a_661_n6069# a_603_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X141 a_287_n2327# a_187_n2415# a_129_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X142 a_n1135_n1109# a_n1235_n1197# a_n1293_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X143 a_n661_n2327# a_n761_n2415# a_n819_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X144 a_n1293_109# a_n1393_21# a_n1451_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X145 a_n503_n3545# a_n603_n3633# a_n661_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X146 a_n819_1327# a_n919_1239# a_n977_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X147 a_287_n3545# a_187_n3633# a_129_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X148 a_n1293_n1109# a_n1393_n1197# a_n1451_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X149 a_n661_1327# a_n761_1239# a_n819_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X150 a_n661_n3545# a_n761_n3633# a_n819_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X151 a_n1135_n2327# a_n1235_n2415# a_n1293_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X152 a_n503_n4763# a_n603_n4851# a_n661_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X153 a_n1451_109# a_n1551_21# a_n1609_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X154 a_1551_n1109# a_1451_n1197# a_1393_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X155 a_n29_n1109# a_n129_n1197# a_n187_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X156 a_n819_2545# a_n919_2457# a_n977_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X157 a_287_n4763# a_187_n4851# a_129_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X158 a_919_1327# a_819_1239# a_761_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X159 a_n1293_n2327# a_n1393_n2415# a_n1451_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X160 a_n661_2545# a_n761_2457# a_n819_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X161 a_n661_n4763# a_n761_n4851# a_n819_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X162 a_n1135_n3545# a_n1235_n3633# a_n1293_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X163 a_n503_n5981# a_n603_n6069# a_n661_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X164 a_n187_n1109# a_n287_n1197# a_n345_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X165 a_n819_3763# a_n919_3675# a_n977_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X166 a_n977_109# a_n1077_21# a_n1135_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X167 a_1551_n2327# a_1451_n2415# a_1393_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X168 a_n29_n2327# a_n129_n2415# a_n187_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X169 a_n187_1327# a_n287_1239# a_n345_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X170 a_761_1327# a_661_1239# a_603_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X171 a_287_n5981# a_187_n6069# a_129_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X172 a_919_2545# a_819_2457# a_761_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X173 a_n1293_n3545# a_n1393_n3633# a_n1451_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X174 a_n661_3763# a_n761_3675# a_n819_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X175 a_n661_n5981# a_n761_n6069# a_n819_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X176 a_n1135_n4763# a_n1235_n4851# a_n1293_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X177 a_n187_n2327# a_n287_n2415# a_n345_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X178 a_n819_4981# a_n919_4893# a_n977_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X179 a_1551_n3545# a_1451_n3633# a_1393_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X180 a_n29_n3545# a_n129_n3633# a_n187_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X181 a_n187_2545# a_n287_2457# a_n345_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X182 a_761_2545# a_661_2457# a_603_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X183 a_n1135_109# a_n1235_21# a_n1293_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X184 a_919_3763# a_819_3675# a_761_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X185 a_n1293_n4763# a_n1393_n4851# a_n1451_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X186 a_n661_4981# a_n761_4893# a_n819_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X187 a_287_1327# a_187_1239# a_129_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X188 a_n1135_n5981# a_n1235_n6069# a_n1293_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X189 a_n187_n3545# a_n287_n3633# a_n345_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X190 a_1551_n4763# a_1451_n4851# a_1393_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X191 a_n29_n4763# a_n129_n4851# a_n187_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X192 a_129_n1109# a_29_n1197# a_n29_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X193 a_761_3763# a_661_3675# a_603_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X194 a_1393_1327# a_1293_1239# a_1235_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X195 a_n187_3763# a_n287_3675# a_n345_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X196 a_n1293_1327# a_n1393_1239# a_n1451_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X197 a_919_4981# a_819_4893# a_761_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X198 a_n1293_n5981# a_n1393_n6069# a_n1451_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X199 a_287_2545# a_187_2457# a_129_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6 a_n108_n250# w_n308_n547# a_50_n250# a_n50_n347#
X0 a_50_n250# a_n50_n347# a_n108_n250# w_n308_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0 a_50_n200# a_n108_n200# a_n50_n288# a_n252_n422#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n252_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_L9TFKV a_n958_n300# a_n900_n388# a_n1092_n522#
+ a_900_n300#
X0 a_900_n300# a_n900_n388# a_n958_n300# a_n1092_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=9
.ends

.subckt sky130_am_ip__ldo_01v8 AVDD VOUT AVSS ENA VREF_EXT SEL_EXT DVDD DVSS
XXM89 AVSS verr AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM56 vbias_p vy AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM78 AVSS AVSS nena ena_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM67 vbias_n vbias_n vbias_n vbias_n AVSS AVSS vbias_n AVSS vbias_n vbias_n vbias_n
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM79 vbias_p vref_int AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM57 vbias_c verr AVDD vy sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM46 vbias_p vx AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM68 AVDD vbias_c vbias_c AVDD sky130_fd_pr__pfet_g5v0d10v5_PC2PN5
Xx1 ENA DVDD DVSS DVSS AVDD AVDD ena_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
XXM58 vbias_c m2_8539_n7649# AVDD vx sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM69 vbias_n vbias_n vbias_c vbias_n AVSS AVSS vbias_c AVSS vbias_c vbias_c vbias_c
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
Xx2 SEL_EXT DVDD DVSS DVSS AVDD AVDD sel_ext_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
XXM59 verr AVSS AVDD vpass sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM48 verr AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXR4 m1_5119_3142# m1_5119_2478# m1_5119_1150# m1_7519_2644# m1_7519_984# m1_7519_1980#
+ m1_5119_2146# m1_5119_3474# m1_7519_1648# m1_5119_1482# m1_7519_2976# m1_5119_2810#
+ vm m1_7519_2976# m1_5119_818# m1_5119_1814# m1_5119_1482# m1_7519_1316# m1_5119_3474#
+ m1_7519_3308# m1_5119_3142# m1_5119_2146# m1_7519_1648# m1_7519_2312# m1_7519_2644#
+ VOUT m1_5119_1150# AVSS m1_5119_2478# m1_7519_1316# m1_5119_2810# m1_7519_3308#
+ m1_7519_2312# m1_5119_818# m1_7519_1980# m1_5119_1814# m1_7519_984# sky130_fd_pr__res_xhigh_po_0p35_QZEXQH
XXR5 m1_5117_n1479# m1_5117_n2475# m1_7517_n4965# m1_5117_n4799# m1_7517_n981# m1_5117_n3803#
+ m1_5117_181# m1_7517_n1977# m1_7517_n3637# m1_7517_n2641# m1_7517_n4633# m1_5117_n815#
+ m1_7517_15# m1_5117_n2475# m1_5117_n5463# m1_5117_n151# m1_5117_n4467# m1_7517_n649#
+ m1_5117_n3471# m1_7517_n2973# m1_5117_n1147# vm m1_7517_n1645# m1_5117_181# m1_5117_n2143#
+ m1_7517_n3969# m1_7517_n4965# m1_5117_n815# m1_5117_n5131# m1_5117_n4135# m1_7517_n1977#
+ m1_5117_n2807# m1_7517_n981# m1_5117_n483# m1_7517_15# m1_7517_n3305# m1_5117_n3139#
+ m1_7517_n4301# m1_7517_n5297# m1_5117_n1479# m1_7517_n1645# m1_7517_n649# m1_7517_n4301#
+ m1_5117_n1811# m1_5117_n2807# m1_7517_n3305# m1_5117_n5463# m1_7517_n5297# m1_5117_n4467#
+ m1_7517_n2641# m1_5117_n151# m1_7517_n2309# m1_7517_n1313# m1_5117_n3471# m1_7517_n317#
+ m1_7517_n4633# m1_5117_n2143# m1_5117_n4799# m1_7517_n3637# AVSS AVSS m1_5117_n1147#
+ m1_5117_n1811# m1_5117_n5131# m1_7517_n1313# m1_5117_n3803# m1_7517_n2309# m1_5117_n483#
+ m1_5117_n4135# m1_7517_n3969# m1_7517_n317# m1_5117_n3139# m1_7517_n2973# sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H
XXR6 AVSS m1_22164_n7435# AVSS m1_22164_n7435# m2_26640_n7437# sky130_fd_pr__res_xhigh_po_0p35_743D3R
XXC1[0] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[1] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[2] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC3 AVSS vref sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM90 nena vdd_start AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM80 vref_int AVSS m1_12626_n9400# m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM70 AVSS vdd_start vbias_n vstart sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM81 vref_int AVSS vref_int m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM71 m1_20910_n7332# vstart vstart AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM60 vbias_p vpass AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM82 vref_int AVSS m1_12626_n9400# AVSS sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM61[0] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[1] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[2] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[3] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[4] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM72 m1_20184_n7334# m1_20910_n7332# m1_20910_n7332# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM83 AVSS AVSS nsel_ext sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM73 AVDD m1_20184_n7334# m1_20184_n7334# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM62 vbias_p AVDD AVDD m1_19028_n7338# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM84 AVDD AVDD nsel_ext sel_ext_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
Xsky130_fd_pr__pfet_g5v0d10v5_KLAZY6_0 ena_3v3 vbias_c AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM63 vbias_c m1_19028_n7338# AVDD vbias_p sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM74 vbias_n vbias_n vstart vbias_n AVSS AVSS vstart AVSS vstart vstart vstart vbias_n
+ AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM85 AVSS vbias_n AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM52 vy m2_6784_n8214# vm AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM53 vx m2_6784_n8214# vref AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM75 AVSS vref vref_int nsel_ext sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM64 vbias_p AVDD AVDD m1_16878_n7330# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM65 vbias_c m1_16878_n7330# AVDD vbias_n sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM87 AVSS vpass AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM54 AVSS vbias_n AVSS m2_6784_n8214# sky130_fd_pr__nfet_g5v0d10v5_L9TFKV
XXM76 AVDD AVDD nena ena_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
XXM66[0] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[1] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[2] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[3] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM55 m2_8539_n7649# AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXM88 ena_3v3 vbias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM77 AVSS VREF_EXT vref sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
.ends

