magic
tech sky130A
magscale 1 2
timestamp 1713187042
<< pwell >>
rect -3106 -1582 3106 1582
<< psubdiff >>
rect -3070 1512 -2974 1546
rect 2974 1512 3070 1546
rect -3070 1450 -3036 1512
rect 3036 1450 3070 1512
rect -3070 -1512 -3036 -1450
rect 3036 -1512 3070 -1450
rect -3070 -1546 -2974 -1512
rect 2974 -1546 3070 -1512
<< psubdiffcont >>
rect -2974 1512 2974 1546
rect -3070 -1450 -3036 1450
rect 3036 -1450 3070 1450
rect -2974 -1546 2974 -1512
<< xpolycontact >>
rect -2940 984 -2870 1416
rect -2940 -1416 -2870 -984
rect -2774 984 -2704 1416
rect -2774 -1416 -2704 -984
rect -2608 984 -2538 1416
rect -2608 -1416 -2538 -984
rect -2442 984 -2372 1416
rect -2442 -1416 -2372 -984
rect -2276 984 -2206 1416
rect -2276 -1416 -2206 -984
rect -2110 984 -2040 1416
rect -2110 -1416 -2040 -984
rect -1944 984 -1874 1416
rect -1944 -1416 -1874 -984
rect -1778 984 -1708 1416
rect -1778 -1416 -1708 -984
rect -1612 984 -1542 1416
rect -1612 -1416 -1542 -984
rect -1446 984 -1376 1416
rect -1446 -1416 -1376 -984
rect -1280 984 -1210 1416
rect -1280 -1416 -1210 -984
rect -1114 984 -1044 1416
rect -1114 -1416 -1044 -984
rect -948 984 -878 1416
rect -948 -1416 -878 -984
rect -782 984 -712 1416
rect -782 -1416 -712 -984
rect -616 984 -546 1416
rect -616 -1416 -546 -984
rect -450 984 -380 1416
rect -450 -1416 -380 -984
rect -284 984 -214 1416
rect -284 -1416 -214 -984
rect -118 984 -48 1416
rect -118 -1416 -48 -984
rect 48 984 118 1416
rect 48 -1416 118 -984
rect 214 984 284 1416
rect 214 -1416 284 -984
rect 380 984 450 1416
rect 380 -1416 450 -984
rect 546 984 616 1416
rect 546 -1416 616 -984
rect 712 984 782 1416
rect 712 -1416 782 -984
rect 878 984 948 1416
rect 878 -1416 948 -984
rect 1044 984 1114 1416
rect 1044 -1416 1114 -984
rect 1210 984 1280 1416
rect 1210 -1416 1280 -984
rect 1376 984 1446 1416
rect 1376 -1416 1446 -984
rect 1542 984 1612 1416
rect 1542 -1416 1612 -984
rect 1708 984 1778 1416
rect 1708 -1416 1778 -984
rect 1874 984 1944 1416
rect 1874 -1416 1944 -984
rect 2040 984 2110 1416
rect 2040 -1416 2110 -984
rect 2206 984 2276 1416
rect 2206 -1416 2276 -984
rect 2372 984 2442 1416
rect 2372 -1416 2442 -984
rect 2538 984 2608 1416
rect 2538 -1416 2608 -984
rect 2704 984 2774 1416
rect 2704 -1416 2774 -984
rect 2870 984 2940 1416
rect 2870 -1416 2940 -984
<< xpolyres >>
rect -2940 -984 -2870 984
rect -2774 -984 -2704 984
rect -2608 -984 -2538 984
rect -2442 -984 -2372 984
rect -2276 -984 -2206 984
rect -2110 -984 -2040 984
rect -1944 -984 -1874 984
rect -1778 -984 -1708 984
rect -1612 -984 -1542 984
rect -1446 -984 -1376 984
rect -1280 -984 -1210 984
rect -1114 -984 -1044 984
rect -948 -984 -878 984
rect -782 -984 -712 984
rect -616 -984 -546 984
rect -450 -984 -380 984
rect -284 -984 -214 984
rect -118 -984 -48 984
rect 48 -984 118 984
rect 214 -984 284 984
rect 380 -984 450 984
rect 546 -984 616 984
rect 712 -984 782 984
rect 878 -984 948 984
rect 1044 -984 1114 984
rect 1210 -984 1280 984
rect 1376 -984 1446 984
rect 1542 -984 1612 984
rect 1708 -984 1778 984
rect 1874 -984 1944 984
rect 2040 -984 2110 984
rect 2206 -984 2276 984
rect 2372 -984 2442 984
rect 2538 -984 2608 984
rect 2704 -984 2774 984
rect 2870 -984 2940 984
<< locali >>
rect -3070 1512 -2974 1546
rect 2974 1512 3070 1546
rect -3070 1450 -3036 1512
rect 3036 1450 3070 1512
rect -3070 -1512 -3036 -1450
rect 3036 -1512 3070 -1450
rect -3070 -1546 -2974 -1512
rect 2974 -1546 3070 -1512
<< viali >>
rect -2924 1001 -2886 1398
rect -2758 1001 -2720 1398
rect -2592 1001 -2554 1398
rect -2426 1001 -2388 1398
rect -2260 1001 -2222 1398
rect -2094 1001 -2056 1398
rect -1928 1001 -1890 1398
rect -1762 1001 -1724 1398
rect -1596 1001 -1558 1398
rect -1430 1001 -1392 1398
rect -1264 1001 -1226 1398
rect -1098 1001 -1060 1398
rect -932 1001 -894 1398
rect -766 1001 -728 1398
rect -600 1001 -562 1398
rect -434 1001 -396 1398
rect -268 1001 -230 1398
rect -102 1001 -64 1398
rect 64 1001 102 1398
rect 230 1001 268 1398
rect 396 1001 434 1398
rect 562 1001 600 1398
rect 728 1001 766 1398
rect 894 1001 932 1398
rect 1060 1001 1098 1398
rect 1226 1001 1264 1398
rect 1392 1001 1430 1398
rect 1558 1001 1596 1398
rect 1724 1001 1762 1398
rect 1890 1001 1928 1398
rect 2056 1001 2094 1398
rect 2222 1001 2260 1398
rect 2388 1001 2426 1398
rect 2554 1001 2592 1398
rect 2720 1001 2758 1398
rect 2886 1001 2924 1398
rect -2924 -1398 -2886 -1001
rect -2758 -1398 -2720 -1001
rect -2592 -1398 -2554 -1001
rect -2426 -1398 -2388 -1001
rect -2260 -1398 -2222 -1001
rect -2094 -1398 -2056 -1001
rect -1928 -1398 -1890 -1001
rect -1762 -1398 -1724 -1001
rect -1596 -1398 -1558 -1001
rect -1430 -1398 -1392 -1001
rect -1264 -1398 -1226 -1001
rect -1098 -1398 -1060 -1001
rect -932 -1398 -894 -1001
rect -766 -1398 -728 -1001
rect -600 -1398 -562 -1001
rect -434 -1398 -396 -1001
rect -268 -1398 -230 -1001
rect -102 -1398 -64 -1001
rect 64 -1398 102 -1001
rect 230 -1398 268 -1001
rect 396 -1398 434 -1001
rect 562 -1398 600 -1001
rect 728 -1398 766 -1001
rect 894 -1398 932 -1001
rect 1060 -1398 1098 -1001
rect 1226 -1398 1264 -1001
rect 1392 -1398 1430 -1001
rect 1558 -1398 1596 -1001
rect 1724 -1398 1762 -1001
rect 1890 -1398 1928 -1001
rect 2056 -1398 2094 -1001
rect 2222 -1398 2260 -1001
rect 2388 -1398 2426 -1001
rect 2554 -1398 2592 -1001
rect 2720 -1398 2758 -1001
rect 2886 -1398 2924 -1001
<< metal1 >>
rect -2930 1398 -2880 1410
rect -2930 1001 -2924 1398
rect -2886 1001 -2880 1398
rect -2930 989 -2880 1001
rect -2764 1398 -2714 1410
rect -2764 1001 -2758 1398
rect -2720 1001 -2714 1398
rect -2764 989 -2714 1001
rect -2598 1398 -2548 1410
rect -2598 1001 -2592 1398
rect -2554 1001 -2548 1398
rect -2598 989 -2548 1001
rect -2432 1398 -2382 1410
rect -2432 1001 -2426 1398
rect -2388 1001 -2382 1398
rect -2432 989 -2382 1001
rect -2266 1398 -2216 1410
rect -2266 1001 -2260 1398
rect -2222 1001 -2216 1398
rect -2266 989 -2216 1001
rect -2100 1398 -2050 1410
rect -2100 1001 -2094 1398
rect -2056 1001 -2050 1398
rect -2100 989 -2050 1001
rect -1934 1398 -1884 1410
rect -1934 1001 -1928 1398
rect -1890 1001 -1884 1398
rect -1934 989 -1884 1001
rect -1768 1398 -1718 1410
rect -1768 1001 -1762 1398
rect -1724 1001 -1718 1398
rect -1768 989 -1718 1001
rect -1602 1398 -1552 1410
rect -1602 1001 -1596 1398
rect -1558 1001 -1552 1398
rect -1602 989 -1552 1001
rect -1436 1398 -1386 1410
rect -1436 1001 -1430 1398
rect -1392 1001 -1386 1398
rect -1436 989 -1386 1001
rect -1270 1398 -1220 1410
rect -1270 1001 -1264 1398
rect -1226 1001 -1220 1398
rect -1270 989 -1220 1001
rect -1104 1398 -1054 1410
rect -1104 1001 -1098 1398
rect -1060 1001 -1054 1398
rect -1104 989 -1054 1001
rect -938 1398 -888 1410
rect -938 1001 -932 1398
rect -894 1001 -888 1398
rect -938 989 -888 1001
rect -772 1398 -722 1410
rect -772 1001 -766 1398
rect -728 1001 -722 1398
rect -772 989 -722 1001
rect -606 1398 -556 1410
rect -606 1001 -600 1398
rect -562 1001 -556 1398
rect -606 989 -556 1001
rect -440 1398 -390 1410
rect -440 1001 -434 1398
rect -396 1001 -390 1398
rect -440 989 -390 1001
rect -274 1398 -224 1410
rect -274 1001 -268 1398
rect -230 1001 -224 1398
rect -274 989 -224 1001
rect -108 1398 -58 1410
rect -108 1001 -102 1398
rect -64 1001 -58 1398
rect -108 989 -58 1001
rect 58 1398 108 1410
rect 58 1001 64 1398
rect 102 1001 108 1398
rect 58 989 108 1001
rect 224 1398 274 1410
rect 224 1001 230 1398
rect 268 1001 274 1398
rect 224 989 274 1001
rect 390 1398 440 1410
rect 390 1001 396 1398
rect 434 1001 440 1398
rect 390 989 440 1001
rect 556 1398 606 1410
rect 556 1001 562 1398
rect 600 1001 606 1398
rect 556 989 606 1001
rect 722 1398 772 1410
rect 722 1001 728 1398
rect 766 1001 772 1398
rect 722 989 772 1001
rect 888 1398 938 1410
rect 888 1001 894 1398
rect 932 1001 938 1398
rect 888 989 938 1001
rect 1054 1398 1104 1410
rect 1054 1001 1060 1398
rect 1098 1001 1104 1398
rect 1054 989 1104 1001
rect 1220 1398 1270 1410
rect 1220 1001 1226 1398
rect 1264 1001 1270 1398
rect 1220 989 1270 1001
rect 1386 1398 1436 1410
rect 1386 1001 1392 1398
rect 1430 1001 1436 1398
rect 1386 989 1436 1001
rect 1552 1398 1602 1410
rect 1552 1001 1558 1398
rect 1596 1001 1602 1398
rect 1552 989 1602 1001
rect 1718 1398 1768 1410
rect 1718 1001 1724 1398
rect 1762 1001 1768 1398
rect 1718 989 1768 1001
rect 1884 1398 1934 1410
rect 1884 1001 1890 1398
rect 1928 1001 1934 1398
rect 1884 989 1934 1001
rect 2050 1398 2100 1410
rect 2050 1001 2056 1398
rect 2094 1001 2100 1398
rect 2050 989 2100 1001
rect 2216 1398 2266 1410
rect 2216 1001 2222 1398
rect 2260 1001 2266 1398
rect 2216 989 2266 1001
rect 2382 1398 2432 1410
rect 2382 1001 2388 1398
rect 2426 1001 2432 1398
rect 2382 989 2432 1001
rect 2548 1398 2598 1410
rect 2548 1001 2554 1398
rect 2592 1001 2598 1398
rect 2548 989 2598 1001
rect 2714 1398 2764 1410
rect 2714 1001 2720 1398
rect 2758 1001 2764 1398
rect 2714 989 2764 1001
rect 2880 1398 2930 1410
rect 2880 1001 2886 1398
rect 2924 1001 2930 1398
rect 2880 989 2930 1001
rect -2930 -1001 -2880 -989
rect -2930 -1398 -2924 -1001
rect -2886 -1398 -2880 -1001
rect -2930 -1410 -2880 -1398
rect -2764 -1001 -2714 -989
rect -2764 -1398 -2758 -1001
rect -2720 -1398 -2714 -1001
rect -2764 -1410 -2714 -1398
rect -2598 -1001 -2548 -989
rect -2598 -1398 -2592 -1001
rect -2554 -1398 -2548 -1001
rect -2598 -1410 -2548 -1398
rect -2432 -1001 -2382 -989
rect -2432 -1398 -2426 -1001
rect -2388 -1398 -2382 -1001
rect -2432 -1410 -2382 -1398
rect -2266 -1001 -2216 -989
rect -2266 -1398 -2260 -1001
rect -2222 -1398 -2216 -1001
rect -2266 -1410 -2216 -1398
rect -2100 -1001 -2050 -989
rect -2100 -1398 -2094 -1001
rect -2056 -1398 -2050 -1001
rect -2100 -1410 -2050 -1398
rect -1934 -1001 -1884 -989
rect -1934 -1398 -1928 -1001
rect -1890 -1398 -1884 -1001
rect -1934 -1410 -1884 -1398
rect -1768 -1001 -1718 -989
rect -1768 -1398 -1762 -1001
rect -1724 -1398 -1718 -1001
rect -1768 -1410 -1718 -1398
rect -1602 -1001 -1552 -989
rect -1602 -1398 -1596 -1001
rect -1558 -1398 -1552 -1001
rect -1602 -1410 -1552 -1398
rect -1436 -1001 -1386 -989
rect -1436 -1398 -1430 -1001
rect -1392 -1398 -1386 -1001
rect -1436 -1410 -1386 -1398
rect -1270 -1001 -1220 -989
rect -1270 -1398 -1264 -1001
rect -1226 -1398 -1220 -1001
rect -1270 -1410 -1220 -1398
rect -1104 -1001 -1054 -989
rect -1104 -1398 -1098 -1001
rect -1060 -1398 -1054 -1001
rect -1104 -1410 -1054 -1398
rect -938 -1001 -888 -989
rect -938 -1398 -932 -1001
rect -894 -1398 -888 -1001
rect -938 -1410 -888 -1398
rect -772 -1001 -722 -989
rect -772 -1398 -766 -1001
rect -728 -1398 -722 -1001
rect -772 -1410 -722 -1398
rect -606 -1001 -556 -989
rect -606 -1398 -600 -1001
rect -562 -1398 -556 -1001
rect -606 -1410 -556 -1398
rect -440 -1001 -390 -989
rect -440 -1398 -434 -1001
rect -396 -1398 -390 -1001
rect -440 -1410 -390 -1398
rect -274 -1001 -224 -989
rect -274 -1398 -268 -1001
rect -230 -1398 -224 -1001
rect -274 -1410 -224 -1398
rect -108 -1001 -58 -989
rect -108 -1398 -102 -1001
rect -64 -1398 -58 -1001
rect -108 -1410 -58 -1398
rect 58 -1001 108 -989
rect 58 -1398 64 -1001
rect 102 -1398 108 -1001
rect 58 -1410 108 -1398
rect 224 -1001 274 -989
rect 224 -1398 230 -1001
rect 268 -1398 274 -1001
rect 224 -1410 274 -1398
rect 390 -1001 440 -989
rect 390 -1398 396 -1001
rect 434 -1398 440 -1001
rect 390 -1410 440 -1398
rect 556 -1001 606 -989
rect 556 -1398 562 -1001
rect 600 -1398 606 -1001
rect 556 -1410 606 -1398
rect 722 -1001 772 -989
rect 722 -1398 728 -1001
rect 766 -1398 772 -1001
rect 722 -1410 772 -1398
rect 888 -1001 938 -989
rect 888 -1398 894 -1001
rect 932 -1398 938 -1001
rect 888 -1410 938 -1398
rect 1054 -1001 1104 -989
rect 1054 -1398 1060 -1001
rect 1098 -1398 1104 -1001
rect 1054 -1410 1104 -1398
rect 1220 -1001 1270 -989
rect 1220 -1398 1226 -1001
rect 1264 -1398 1270 -1001
rect 1220 -1410 1270 -1398
rect 1386 -1001 1436 -989
rect 1386 -1398 1392 -1001
rect 1430 -1398 1436 -1001
rect 1386 -1410 1436 -1398
rect 1552 -1001 1602 -989
rect 1552 -1398 1558 -1001
rect 1596 -1398 1602 -1001
rect 1552 -1410 1602 -1398
rect 1718 -1001 1768 -989
rect 1718 -1398 1724 -1001
rect 1762 -1398 1768 -1001
rect 1718 -1410 1768 -1398
rect 1884 -1001 1934 -989
rect 1884 -1398 1890 -1001
rect 1928 -1398 1934 -1001
rect 1884 -1410 1934 -1398
rect 2050 -1001 2100 -989
rect 2050 -1398 2056 -1001
rect 2094 -1398 2100 -1001
rect 2050 -1410 2100 -1398
rect 2216 -1001 2266 -989
rect 2216 -1398 2222 -1001
rect 2260 -1398 2266 -1001
rect 2216 -1410 2266 -1398
rect 2382 -1001 2432 -989
rect 2382 -1398 2388 -1001
rect 2426 -1398 2432 -1001
rect 2382 -1410 2432 -1398
rect 2548 -1001 2598 -989
rect 2548 -1398 2554 -1001
rect 2592 -1398 2598 -1001
rect 2548 -1410 2598 -1398
rect 2714 -1001 2764 -989
rect 2714 -1398 2720 -1001
rect 2758 -1398 2764 -1001
rect 2714 -1410 2764 -1398
rect 2880 -1001 2930 -989
rect 2880 -1398 2886 -1001
rect 2924 -1398 2930 -1001
rect 2880 -1410 2930 -1398
<< properties >>
string FIXED_BBOX -3053 -1529 3053 1529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10.0 m 1 nx 36 wmin 0.350 lmin 0.50 rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
