magic
tech sky130A
timestamp 1713186496
<< pwell >>
rect -214 -179 214 179
<< mvnmos >>
rect -100 -50 100 50
<< mvndiff >>
rect -129 44 -100 50
rect -129 -44 -123 44
rect -106 -44 -100 44
rect -129 -50 -100 -44
rect 100 44 129 50
rect 100 -44 106 44
rect 123 -44 129 44
rect 100 -50 129 -44
<< mvndiffc >>
rect -123 -44 -106 44
rect 106 -44 123 44
<< mvpsubdiff >>
rect -196 155 196 161
rect -196 138 -142 155
rect 142 138 196 155
rect -196 132 196 138
rect -196 107 -167 132
rect -196 -107 -190 107
rect -173 -107 -167 107
rect 167 107 196 132
rect -196 -132 -167 -107
rect 167 -107 173 107
rect 190 -107 196 107
rect 167 -132 196 -107
rect -196 -138 196 -132
rect -196 -155 -142 -138
rect 142 -155 196 -138
rect -196 -161 196 -155
<< mvpsubdiffcont >>
rect -142 138 142 155
rect -190 -107 -173 107
rect 173 -107 190 107
rect -142 -155 142 -138
<< poly >>
rect -100 86 100 94
rect -100 69 -92 86
rect 92 69 100 86
rect -100 50 100 69
rect -100 -69 100 -50
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -100 -94 100 -86
<< polycont >>
rect -92 69 92 86
rect -92 -86 92 -69
<< locali >>
rect -190 138 -142 155
rect 142 138 190 155
rect -190 107 -173 138
rect 173 107 190 138
rect -100 69 -92 86
rect 92 69 100 86
rect -123 44 -106 52
rect -123 -52 -106 -44
rect 106 44 123 52
rect 106 -52 123 -44
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -190 -138 -173 -107
rect 173 -138 190 -107
rect -190 -155 -142 -138
rect 142 -155 190 -138
<< viali >>
rect -92 69 92 86
rect -123 -44 -106 44
rect 106 -44 123 44
rect -92 -86 92 -69
<< metal1 >>
rect -98 86 98 89
rect -98 69 -92 86
rect 92 69 98 86
rect -98 66 98 69
rect -126 44 -103 50
rect -126 -44 -123 44
rect -106 -44 -103 44
rect -126 -50 -103 -44
rect 103 44 126 50
rect 103 -44 106 44
rect 123 -44 126 44
rect 103 -50 126 -44
rect -98 -69 98 -66
rect -98 -86 -92 -69
rect 92 -86 98 -69
rect -98 -89 98 -86
<< properties >>
string FIXED_BBOX -181 -146 181 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
