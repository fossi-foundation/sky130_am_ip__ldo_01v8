magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< metal3 >>
rect -536 362 536 390
rect -536 -362 452 362
rect 516 -362 536 362
rect -536 -390 536 -362
<< via3 >>
rect 452 -362 516 362
<< mimcap >>
rect -496 310 204 350
rect -496 -310 -456 310
rect 164 -310 204 310
rect -496 -350 204 -310
<< mimcapcontact >>
rect -456 -310 164 310
<< metal4 >>
rect 436 362 532 378
rect -457 310 165 311
rect -457 -310 -456 310
rect 164 -310 165 310
rect -457 -311 165 -310
rect 436 -362 452 362
rect 516 -362 532 362
rect 436 -378 532 -362
<< properties >>
string FIXED_BBOX -536 -390 244 390
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.5 l 3.5 val 27.16 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
