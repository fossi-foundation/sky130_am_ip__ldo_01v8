magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -1258 -615 1258 615
<< mvpmos >>
rect -1000 118 1000 318
rect -1000 -318 1000 -118
<< mvpdiff >>
rect -1058 306 -1000 318
rect -1058 130 -1046 306
rect -1012 130 -1000 306
rect -1058 118 -1000 130
rect 1000 306 1058 318
rect 1000 130 1012 306
rect 1046 130 1058 306
rect 1000 118 1058 130
rect -1058 -130 -1000 -118
rect -1058 -306 -1046 -130
rect -1012 -306 -1000 -130
rect -1058 -318 -1000 -306
rect 1000 -130 1058 -118
rect 1000 -306 1012 -130
rect 1046 -306 1058 -130
rect 1000 -318 1058 -306
<< mvpdiffc >>
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
<< mvnsubdiff >>
rect -1192 537 1192 549
rect -1192 503 -1084 537
rect 1084 503 1192 537
rect -1192 491 1192 503
rect -1192 441 -1134 491
rect -1192 -441 -1180 441
rect -1146 -441 -1134 441
rect 1134 441 1192 491
rect -1192 -491 -1134 -441
rect 1134 -441 1146 441
rect 1180 -441 1192 441
rect 1134 -491 1192 -441
rect -1192 -503 1192 -491
rect -1192 -537 -1084 -503
rect 1084 -537 1192 -503
rect -1192 -549 1192 -537
<< mvnsubdiffcont >>
rect -1084 503 1084 537
rect -1180 -441 -1146 441
rect 1146 -441 1180 441
rect -1084 -537 1084 -503
<< poly >>
rect -1000 399 1000 415
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1000 318 1000 365
rect -1000 71 1000 118
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -118 1000 -71
rect -1000 -365 1000 -318
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1000 -415 1000 -399
<< polycont >>
rect -984 365 984 399
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -399 984 -365
<< locali >>
rect -1180 503 -1084 537
rect 1084 503 1180 537
rect -1180 441 -1146 503
rect 1146 441 1180 503
rect -1000 365 -984 399
rect 984 365 1000 399
rect -1046 306 -1012 322
rect -1046 114 -1012 130
rect 1012 306 1046 322
rect 1012 114 1046 130
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -130 -1012 -114
rect -1046 -322 -1012 -306
rect 1012 -130 1046 -114
rect 1012 -322 1046 -306
rect -1000 -399 -984 -365
rect 984 -399 1000 -365
rect -1180 -503 -1146 -441
rect 1146 -503 1180 -441
rect -1180 -537 -1084 -503
rect 1084 -537 1180 -503
<< viali >>
rect -984 365 984 399
rect -1046 130 -1012 306
rect 1012 130 1046 306
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -306 -1012 -130
rect 1012 -306 1046 -130
rect -984 -399 984 -365
<< metal1 >>
rect -996 399 996 405
rect -996 365 -984 399
rect 984 365 996 399
rect -996 359 996 365
rect -1052 306 -1006 318
rect -1052 130 -1046 306
rect -1012 130 -1006 306
rect -1052 118 -1006 130
rect 1006 306 1052 318
rect 1006 130 1012 306
rect 1046 130 1052 306
rect 1006 118 1052 130
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -130 -1006 -118
rect -1052 -306 -1046 -130
rect -1012 -306 -1006 -130
rect -1052 -318 -1006 -306
rect 1006 -130 1052 -118
rect 1006 -306 1012 -130
rect 1046 -306 1052 -130
rect 1006 -318 1052 -306
rect -996 -365 996 -359
rect -996 -399 -984 -365
rect 984 -399 996 -365
rect -996 -405 996 -399
<< properties >>
string FIXED_BBOX -1163 -520 1163 520
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
