magic
tech sky130A
magscale 1 2
timestamp 1717294357
<< nwell >>
rect -458 -397 458 397
<< mvpmos >>
rect -200 -100 200 100
<< mvpdiff >>
rect -258 88 -200 100
rect -258 -88 -246 88
rect -212 -88 -200 88
rect -258 -100 -200 -88
rect 200 88 258 100
rect 200 -88 212 88
rect 246 -88 258 88
rect 200 -100 258 -88
<< mvpdiffc >>
rect -246 -88 -212 88
rect 212 -88 246 88
<< mvnsubdiff >>
rect -392 319 392 331
rect -392 285 -284 319
rect 284 285 392 319
rect -392 273 392 285
rect -392 223 -334 273
rect -392 -223 -380 223
rect -346 -223 -334 223
rect 334 223 392 273
rect -392 -273 -334 -223
rect 334 -223 346 223
rect 380 -223 392 223
rect 334 -273 392 -223
rect -392 -285 392 -273
rect -392 -319 -284 -285
rect 284 -319 392 -285
rect -392 -331 392 -319
<< mvnsubdiffcont >>
rect -284 285 284 319
rect -380 -223 -346 223
rect 346 -223 380 223
rect -284 -319 284 -285
<< poly >>
rect -200 181 200 197
rect -200 147 -184 181
rect 184 147 200 181
rect -200 100 200 147
rect -200 -147 200 -100
rect -200 -181 -184 -147
rect 184 -181 200 -147
rect -200 -197 200 -181
<< polycont >>
rect -184 147 184 181
rect -184 -181 184 -147
<< locali >>
rect -380 285 -284 319
rect 284 285 380 319
rect -380 223 -346 285
rect 346 223 380 285
rect -200 147 -184 181
rect 184 147 200 181
rect -246 88 -212 104
rect -246 -104 -212 -88
rect 212 88 246 104
rect 212 -104 246 -88
rect -200 -181 -184 -147
rect 184 -181 200 -147
rect -380 -285 -346 -223
rect 346 -285 380 -223
rect -380 -319 -284 -285
rect 284 -319 380 -285
<< viali >>
rect -184 147 184 181
rect -246 -88 -212 88
rect 212 -88 246 88
rect -184 -181 184 -147
<< metal1 >>
rect -196 181 196 187
rect -196 147 -184 181
rect 184 147 196 181
rect -196 141 196 147
rect -252 88 -206 100
rect -252 -88 -246 88
rect -212 -88 -206 88
rect -252 -100 -206 -88
rect 206 88 252 100
rect 206 -88 212 88
rect 246 -88 252 88
rect 206 -100 252 -88
rect -196 -147 196 -141
rect -196 -181 -184 -147
rect 184 -181 196 -147
rect -196 -187 196 -181
<< properties >>
string FIXED_BBOX -363 -302 363 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
