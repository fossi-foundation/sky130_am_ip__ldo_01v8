magic
tech sky130A
magscale 1 2
timestamp 1717253844
<< pwell >>
rect -278 -609149 278 609149
<< mvnmos >>
rect -50 607891 50 608891
rect -50 606673 50 607673
rect -50 605455 50 606455
rect -50 604237 50 605237
rect -50 603019 50 604019
rect -50 601801 50 602801
rect -50 600583 50 601583
rect -50 599365 50 600365
rect -50 598147 50 599147
rect -50 596929 50 597929
rect -50 595711 50 596711
rect -50 594493 50 595493
rect -50 593275 50 594275
rect -50 592057 50 593057
rect -50 590839 50 591839
rect -50 589621 50 590621
rect -50 588403 50 589403
rect -50 587185 50 588185
rect -50 585967 50 586967
rect -50 584749 50 585749
rect -50 583531 50 584531
rect -50 582313 50 583313
rect -50 581095 50 582095
rect -50 579877 50 580877
rect -50 578659 50 579659
rect -50 577441 50 578441
rect -50 576223 50 577223
rect -50 575005 50 576005
rect -50 573787 50 574787
rect -50 572569 50 573569
rect -50 571351 50 572351
rect -50 570133 50 571133
rect -50 568915 50 569915
rect -50 567697 50 568697
rect -50 566479 50 567479
rect -50 565261 50 566261
rect -50 564043 50 565043
rect -50 562825 50 563825
rect -50 561607 50 562607
rect -50 560389 50 561389
rect -50 559171 50 560171
rect -50 557953 50 558953
rect -50 556735 50 557735
rect -50 555517 50 556517
rect -50 554299 50 555299
rect -50 553081 50 554081
rect -50 551863 50 552863
rect -50 550645 50 551645
rect -50 549427 50 550427
rect -50 548209 50 549209
rect -50 546991 50 547991
rect -50 545773 50 546773
rect -50 544555 50 545555
rect -50 543337 50 544337
rect -50 542119 50 543119
rect -50 540901 50 541901
rect -50 539683 50 540683
rect -50 538465 50 539465
rect -50 537247 50 538247
rect -50 536029 50 537029
rect -50 534811 50 535811
rect -50 533593 50 534593
rect -50 532375 50 533375
rect -50 531157 50 532157
rect -50 529939 50 530939
rect -50 528721 50 529721
rect -50 527503 50 528503
rect -50 526285 50 527285
rect -50 525067 50 526067
rect -50 523849 50 524849
rect -50 522631 50 523631
rect -50 521413 50 522413
rect -50 520195 50 521195
rect -50 518977 50 519977
rect -50 517759 50 518759
rect -50 516541 50 517541
rect -50 515323 50 516323
rect -50 514105 50 515105
rect -50 512887 50 513887
rect -50 511669 50 512669
rect -50 510451 50 511451
rect -50 509233 50 510233
rect -50 508015 50 509015
rect -50 506797 50 507797
rect -50 505579 50 506579
rect -50 504361 50 505361
rect -50 503143 50 504143
rect -50 501925 50 502925
rect -50 500707 50 501707
rect -50 499489 50 500489
rect -50 498271 50 499271
rect -50 497053 50 498053
rect -50 495835 50 496835
rect -50 494617 50 495617
rect -50 493399 50 494399
rect -50 492181 50 493181
rect -50 490963 50 491963
rect -50 489745 50 490745
rect -50 488527 50 489527
rect -50 487309 50 488309
rect -50 486091 50 487091
rect -50 484873 50 485873
rect -50 483655 50 484655
rect -50 482437 50 483437
rect -50 481219 50 482219
rect -50 480001 50 481001
rect -50 478783 50 479783
rect -50 477565 50 478565
rect -50 476347 50 477347
rect -50 475129 50 476129
rect -50 473911 50 474911
rect -50 472693 50 473693
rect -50 471475 50 472475
rect -50 470257 50 471257
rect -50 469039 50 470039
rect -50 467821 50 468821
rect -50 466603 50 467603
rect -50 465385 50 466385
rect -50 464167 50 465167
rect -50 462949 50 463949
rect -50 461731 50 462731
rect -50 460513 50 461513
rect -50 459295 50 460295
rect -50 458077 50 459077
rect -50 456859 50 457859
rect -50 455641 50 456641
rect -50 454423 50 455423
rect -50 453205 50 454205
rect -50 451987 50 452987
rect -50 450769 50 451769
rect -50 449551 50 450551
rect -50 448333 50 449333
rect -50 447115 50 448115
rect -50 445897 50 446897
rect -50 444679 50 445679
rect -50 443461 50 444461
rect -50 442243 50 443243
rect -50 441025 50 442025
rect -50 439807 50 440807
rect -50 438589 50 439589
rect -50 437371 50 438371
rect -50 436153 50 437153
rect -50 434935 50 435935
rect -50 433717 50 434717
rect -50 432499 50 433499
rect -50 431281 50 432281
rect -50 430063 50 431063
rect -50 428845 50 429845
rect -50 427627 50 428627
rect -50 426409 50 427409
rect -50 425191 50 426191
rect -50 423973 50 424973
rect -50 422755 50 423755
rect -50 421537 50 422537
rect -50 420319 50 421319
rect -50 419101 50 420101
rect -50 417883 50 418883
rect -50 416665 50 417665
rect -50 415447 50 416447
rect -50 414229 50 415229
rect -50 413011 50 414011
rect -50 411793 50 412793
rect -50 410575 50 411575
rect -50 409357 50 410357
rect -50 408139 50 409139
rect -50 406921 50 407921
rect -50 405703 50 406703
rect -50 404485 50 405485
rect -50 403267 50 404267
rect -50 402049 50 403049
rect -50 400831 50 401831
rect -50 399613 50 400613
rect -50 398395 50 399395
rect -50 397177 50 398177
rect -50 395959 50 396959
rect -50 394741 50 395741
rect -50 393523 50 394523
rect -50 392305 50 393305
rect -50 391087 50 392087
rect -50 389869 50 390869
rect -50 388651 50 389651
rect -50 387433 50 388433
rect -50 386215 50 387215
rect -50 384997 50 385997
rect -50 383779 50 384779
rect -50 382561 50 383561
rect -50 381343 50 382343
rect -50 380125 50 381125
rect -50 378907 50 379907
rect -50 377689 50 378689
rect -50 376471 50 377471
rect -50 375253 50 376253
rect -50 374035 50 375035
rect -50 372817 50 373817
rect -50 371599 50 372599
rect -50 370381 50 371381
rect -50 369163 50 370163
rect -50 367945 50 368945
rect -50 366727 50 367727
rect -50 365509 50 366509
rect -50 364291 50 365291
rect -50 363073 50 364073
rect -50 361855 50 362855
rect -50 360637 50 361637
rect -50 359419 50 360419
rect -50 358201 50 359201
rect -50 356983 50 357983
rect -50 355765 50 356765
rect -50 354547 50 355547
rect -50 353329 50 354329
rect -50 352111 50 353111
rect -50 350893 50 351893
rect -50 349675 50 350675
rect -50 348457 50 349457
rect -50 347239 50 348239
rect -50 346021 50 347021
rect -50 344803 50 345803
rect -50 343585 50 344585
rect -50 342367 50 343367
rect -50 341149 50 342149
rect -50 339931 50 340931
rect -50 338713 50 339713
rect -50 337495 50 338495
rect -50 336277 50 337277
rect -50 335059 50 336059
rect -50 333841 50 334841
rect -50 332623 50 333623
rect -50 331405 50 332405
rect -50 330187 50 331187
rect -50 328969 50 329969
rect -50 327751 50 328751
rect -50 326533 50 327533
rect -50 325315 50 326315
rect -50 324097 50 325097
rect -50 322879 50 323879
rect -50 321661 50 322661
rect -50 320443 50 321443
rect -50 319225 50 320225
rect -50 318007 50 319007
rect -50 316789 50 317789
rect -50 315571 50 316571
rect -50 314353 50 315353
rect -50 313135 50 314135
rect -50 311917 50 312917
rect -50 310699 50 311699
rect -50 309481 50 310481
rect -50 308263 50 309263
rect -50 307045 50 308045
rect -50 305827 50 306827
rect -50 304609 50 305609
rect -50 303391 50 304391
rect -50 302173 50 303173
rect -50 300955 50 301955
rect -50 299737 50 300737
rect -50 298519 50 299519
rect -50 297301 50 298301
rect -50 296083 50 297083
rect -50 294865 50 295865
rect -50 293647 50 294647
rect -50 292429 50 293429
rect -50 291211 50 292211
rect -50 289993 50 290993
rect -50 288775 50 289775
rect -50 287557 50 288557
rect -50 286339 50 287339
rect -50 285121 50 286121
rect -50 283903 50 284903
rect -50 282685 50 283685
rect -50 281467 50 282467
rect -50 280249 50 281249
rect -50 279031 50 280031
rect -50 277813 50 278813
rect -50 276595 50 277595
rect -50 275377 50 276377
rect -50 274159 50 275159
rect -50 272941 50 273941
rect -50 271723 50 272723
rect -50 270505 50 271505
rect -50 269287 50 270287
rect -50 268069 50 269069
rect -50 266851 50 267851
rect -50 265633 50 266633
rect -50 264415 50 265415
rect -50 263197 50 264197
rect -50 261979 50 262979
rect -50 260761 50 261761
rect -50 259543 50 260543
rect -50 258325 50 259325
rect -50 257107 50 258107
rect -50 255889 50 256889
rect -50 254671 50 255671
rect -50 253453 50 254453
rect -50 252235 50 253235
rect -50 251017 50 252017
rect -50 249799 50 250799
rect -50 248581 50 249581
rect -50 247363 50 248363
rect -50 246145 50 247145
rect -50 244927 50 245927
rect -50 243709 50 244709
rect -50 242491 50 243491
rect -50 241273 50 242273
rect -50 240055 50 241055
rect -50 238837 50 239837
rect -50 237619 50 238619
rect -50 236401 50 237401
rect -50 235183 50 236183
rect -50 233965 50 234965
rect -50 232747 50 233747
rect -50 231529 50 232529
rect -50 230311 50 231311
rect -50 229093 50 230093
rect -50 227875 50 228875
rect -50 226657 50 227657
rect -50 225439 50 226439
rect -50 224221 50 225221
rect -50 223003 50 224003
rect -50 221785 50 222785
rect -50 220567 50 221567
rect -50 219349 50 220349
rect -50 218131 50 219131
rect -50 216913 50 217913
rect -50 215695 50 216695
rect -50 214477 50 215477
rect -50 213259 50 214259
rect -50 212041 50 213041
rect -50 210823 50 211823
rect -50 209605 50 210605
rect -50 208387 50 209387
rect -50 207169 50 208169
rect -50 205951 50 206951
rect -50 204733 50 205733
rect -50 203515 50 204515
rect -50 202297 50 203297
rect -50 201079 50 202079
rect -50 199861 50 200861
rect -50 198643 50 199643
rect -50 197425 50 198425
rect -50 196207 50 197207
rect -50 194989 50 195989
rect -50 193771 50 194771
rect -50 192553 50 193553
rect -50 191335 50 192335
rect -50 190117 50 191117
rect -50 188899 50 189899
rect -50 187681 50 188681
rect -50 186463 50 187463
rect -50 185245 50 186245
rect -50 184027 50 185027
rect -50 182809 50 183809
rect -50 181591 50 182591
rect -50 180373 50 181373
rect -50 179155 50 180155
rect -50 177937 50 178937
rect -50 176719 50 177719
rect -50 175501 50 176501
rect -50 174283 50 175283
rect -50 173065 50 174065
rect -50 171847 50 172847
rect -50 170629 50 171629
rect -50 169411 50 170411
rect -50 168193 50 169193
rect -50 166975 50 167975
rect -50 165757 50 166757
rect -50 164539 50 165539
rect -50 163321 50 164321
rect -50 162103 50 163103
rect -50 160885 50 161885
rect -50 159667 50 160667
rect -50 158449 50 159449
rect -50 157231 50 158231
rect -50 156013 50 157013
rect -50 154795 50 155795
rect -50 153577 50 154577
rect -50 152359 50 153359
rect -50 151141 50 152141
rect -50 149923 50 150923
rect -50 148705 50 149705
rect -50 147487 50 148487
rect -50 146269 50 147269
rect -50 145051 50 146051
rect -50 143833 50 144833
rect -50 142615 50 143615
rect -50 141397 50 142397
rect -50 140179 50 141179
rect -50 138961 50 139961
rect -50 137743 50 138743
rect -50 136525 50 137525
rect -50 135307 50 136307
rect -50 134089 50 135089
rect -50 132871 50 133871
rect -50 131653 50 132653
rect -50 130435 50 131435
rect -50 129217 50 130217
rect -50 127999 50 128999
rect -50 126781 50 127781
rect -50 125563 50 126563
rect -50 124345 50 125345
rect -50 123127 50 124127
rect -50 121909 50 122909
rect -50 120691 50 121691
rect -50 119473 50 120473
rect -50 118255 50 119255
rect -50 117037 50 118037
rect -50 115819 50 116819
rect -50 114601 50 115601
rect -50 113383 50 114383
rect -50 112165 50 113165
rect -50 110947 50 111947
rect -50 109729 50 110729
rect -50 108511 50 109511
rect -50 107293 50 108293
rect -50 106075 50 107075
rect -50 104857 50 105857
rect -50 103639 50 104639
rect -50 102421 50 103421
rect -50 101203 50 102203
rect -50 99985 50 100985
rect -50 98767 50 99767
rect -50 97549 50 98549
rect -50 96331 50 97331
rect -50 95113 50 96113
rect -50 93895 50 94895
rect -50 92677 50 93677
rect -50 91459 50 92459
rect -50 90241 50 91241
rect -50 89023 50 90023
rect -50 87805 50 88805
rect -50 86587 50 87587
rect -50 85369 50 86369
rect -50 84151 50 85151
rect -50 82933 50 83933
rect -50 81715 50 82715
rect -50 80497 50 81497
rect -50 79279 50 80279
rect -50 78061 50 79061
rect -50 76843 50 77843
rect -50 75625 50 76625
rect -50 74407 50 75407
rect -50 73189 50 74189
rect -50 71971 50 72971
rect -50 70753 50 71753
rect -50 69535 50 70535
rect -50 68317 50 69317
rect -50 67099 50 68099
rect -50 65881 50 66881
rect -50 64663 50 65663
rect -50 63445 50 64445
rect -50 62227 50 63227
rect -50 61009 50 62009
rect -50 59791 50 60791
rect -50 58573 50 59573
rect -50 57355 50 58355
rect -50 56137 50 57137
rect -50 54919 50 55919
rect -50 53701 50 54701
rect -50 52483 50 53483
rect -50 51265 50 52265
rect -50 50047 50 51047
rect -50 48829 50 49829
rect -50 47611 50 48611
rect -50 46393 50 47393
rect -50 45175 50 46175
rect -50 43957 50 44957
rect -50 42739 50 43739
rect -50 41521 50 42521
rect -50 40303 50 41303
rect -50 39085 50 40085
rect -50 37867 50 38867
rect -50 36649 50 37649
rect -50 35431 50 36431
rect -50 34213 50 35213
rect -50 32995 50 33995
rect -50 31777 50 32777
rect -50 30559 50 31559
rect -50 29341 50 30341
rect -50 28123 50 29123
rect -50 26905 50 27905
rect -50 25687 50 26687
rect -50 24469 50 25469
rect -50 23251 50 24251
rect -50 22033 50 23033
rect -50 20815 50 21815
rect -50 19597 50 20597
rect -50 18379 50 19379
rect -50 17161 50 18161
rect -50 15943 50 16943
rect -50 14725 50 15725
rect -50 13507 50 14507
rect -50 12289 50 13289
rect -50 11071 50 12071
rect -50 9853 50 10853
rect -50 8635 50 9635
rect -50 7417 50 8417
rect -50 6199 50 7199
rect -50 4981 50 5981
rect -50 3763 50 4763
rect -50 2545 50 3545
rect -50 1327 50 2327
rect -50 109 50 1109
rect -50 -1109 50 -109
rect -50 -2327 50 -1327
rect -50 -3545 50 -2545
rect -50 -4763 50 -3763
rect -50 -5981 50 -4981
rect -50 -7199 50 -6199
rect -50 -8417 50 -7417
rect -50 -9635 50 -8635
rect -50 -10853 50 -9853
rect -50 -12071 50 -11071
rect -50 -13289 50 -12289
rect -50 -14507 50 -13507
rect -50 -15725 50 -14725
rect -50 -16943 50 -15943
rect -50 -18161 50 -17161
rect -50 -19379 50 -18379
rect -50 -20597 50 -19597
rect -50 -21815 50 -20815
rect -50 -23033 50 -22033
rect -50 -24251 50 -23251
rect -50 -25469 50 -24469
rect -50 -26687 50 -25687
rect -50 -27905 50 -26905
rect -50 -29123 50 -28123
rect -50 -30341 50 -29341
rect -50 -31559 50 -30559
rect -50 -32777 50 -31777
rect -50 -33995 50 -32995
rect -50 -35213 50 -34213
rect -50 -36431 50 -35431
rect -50 -37649 50 -36649
rect -50 -38867 50 -37867
rect -50 -40085 50 -39085
rect -50 -41303 50 -40303
rect -50 -42521 50 -41521
rect -50 -43739 50 -42739
rect -50 -44957 50 -43957
rect -50 -46175 50 -45175
rect -50 -47393 50 -46393
rect -50 -48611 50 -47611
rect -50 -49829 50 -48829
rect -50 -51047 50 -50047
rect -50 -52265 50 -51265
rect -50 -53483 50 -52483
rect -50 -54701 50 -53701
rect -50 -55919 50 -54919
rect -50 -57137 50 -56137
rect -50 -58355 50 -57355
rect -50 -59573 50 -58573
rect -50 -60791 50 -59791
rect -50 -62009 50 -61009
rect -50 -63227 50 -62227
rect -50 -64445 50 -63445
rect -50 -65663 50 -64663
rect -50 -66881 50 -65881
rect -50 -68099 50 -67099
rect -50 -69317 50 -68317
rect -50 -70535 50 -69535
rect -50 -71753 50 -70753
rect -50 -72971 50 -71971
rect -50 -74189 50 -73189
rect -50 -75407 50 -74407
rect -50 -76625 50 -75625
rect -50 -77843 50 -76843
rect -50 -79061 50 -78061
rect -50 -80279 50 -79279
rect -50 -81497 50 -80497
rect -50 -82715 50 -81715
rect -50 -83933 50 -82933
rect -50 -85151 50 -84151
rect -50 -86369 50 -85369
rect -50 -87587 50 -86587
rect -50 -88805 50 -87805
rect -50 -90023 50 -89023
rect -50 -91241 50 -90241
rect -50 -92459 50 -91459
rect -50 -93677 50 -92677
rect -50 -94895 50 -93895
rect -50 -96113 50 -95113
rect -50 -97331 50 -96331
rect -50 -98549 50 -97549
rect -50 -99767 50 -98767
rect -50 -100985 50 -99985
rect -50 -102203 50 -101203
rect -50 -103421 50 -102421
rect -50 -104639 50 -103639
rect -50 -105857 50 -104857
rect -50 -107075 50 -106075
rect -50 -108293 50 -107293
rect -50 -109511 50 -108511
rect -50 -110729 50 -109729
rect -50 -111947 50 -110947
rect -50 -113165 50 -112165
rect -50 -114383 50 -113383
rect -50 -115601 50 -114601
rect -50 -116819 50 -115819
rect -50 -118037 50 -117037
rect -50 -119255 50 -118255
rect -50 -120473 50 -119473
rect -50 -121691 50 -120691
rect -50 -122909 50 -121909
rect -50 -124127 50 -123127
rect -50 -125345 50 -124345
rect -50 -126563 50 -125563
rect -50 -127781 50 -126781
rect -50 -128999 50 -127999
rect -50 -130217 50 -129217
rect -50 -131435 50 -130435
rect -50 -132653 50 -131653
rect -50 -133871 50 -132871
rect -50 -135089 50 -134089
rect -50 -136307 50 -135307
rect -50 -137525 50 -136525
rect -50 -138743 50 -137743
rect -50 -139961 50 -138961
rect -50 -141179 50 -140179
rect -50 -142397 50 -141397
rect -50 -143615 50 -142615
rect -50 -144833 50 -143833
rect -50 -146051 50 -145051
rect -50 -147269 50 -146269
rect -50 -148487 50 -147487
rect -50 -149705 50 -148705
rect -50 -150923 50 -149923
rect -50 -152141 50 -151141
rect -50 -153359 50 -152359
rect -50 -154577 50 -153577
rect -50 -155795 50 -154795
rect -50 -157013 50 -156013
rect -50 -158231 50 -157231
rect -50 -159449 50 -158449
rect -50 -160667 50 -159667
rect -50 -161885 50 -160885
rect -50 -163103 50 -162103
rect -50 -164321 50 -163321
rect -50 -165539 50 -164539
rect -50 -166757 50 -165757
rect -50 -167975 50 -166975
rect -50 -169193 50 -168193
rect -50 -170411 50 -169411
rect -50 -171629 50 -170629
rect -50 -172847 50 -171847
rect -50 -174065 50 -173065
rect -50 -175283 50 -174283
rect -50 -176501 50 -175501
rect -50 -177719 50 -176719
rect -50 -178937 50 -177937
rect -50 -180155 50 -179155
rect -50 -181373 50 -180373
rect -50 -182591 50 -181591
rect -50 -183809 50 -182809
rect -50 -185027 50 -184027
rect -50 -186245 50 -185245
rect -50 -187463 50 -186463
rect -50 -188681 50 -187681
rect -50 -189899 50 -188899
rect -50 -191117 50 -190117
rect -50 -192335 50 -191335
rect -50 -193553 50 -192553
rect -50 -194771 50 -193771
rect -50 -195989 50 -194989
rect -50 -197207 50 -196207
rect -50 -198425 50 -197425
rect -50 -199643 50 -198643
rect -50 -200861 50 -199861
rect -50 -202079 50 -201079
rect -50 -203297 50 -202297
rect -50 -204515 50 -203515
rect -50 -205733 50 -204733
rect -50 -206951 50 -205951
rect -50 -208169 50 -207169
rect -50 -209387 50 -208387
rect -50 -210605 50 -209605
rect -50 -211823 50 -210823
rect -50 -213041 50 -212041
rect -50 -214259 50 -213259
rect -50 -215477 50 -214477
rect -50 -216695 50 -215695
rect -50 -217913 50 -216913
rect -50 -219131 50 -218131
rect -50 -220349 50 -219349
rect -50 -221567 50 -220567
rect -50 -222785 50 -221785
rect -50 -224003 50 -223003
rect -50 -225221 50 -224221
rect -50 -226439 50 -225439
rect -50 -227657 50 -226657
rect -50 -228875 50 -227875
rect -50 -230093 50 -229093
rect -50 -231311 50 -230311
rect -50 -232529 50 -231529
rect -50 -233747 50 -232747
rect -50 -234965 50 -233965
rect -50 -236183 50 -235183
rect -50 -237401 50 -236401
rect -50 -238619 50 -237619
rect -50 -239837 50 -238837
rect -50 -241055 50 -240055
rect -50 -242273 50 -241273
rect -50 -243491 50 -242491
rect -50 -244709 50 -243709
rect -50 -245927 50 -244927
rect -50 -247145 50 -246145
rect -50 -248363 50 -247363
rect -50 -249581 50 -248581
rect -50 -250799 50 -249799
rect -50 -252017 50 -251017
rect -50 -253235 50 -252235
rect -50 -254453 50 -253453
rect -50 -255671 50 -254671
rect -50 -256889 50 -255889
rect -50 -258107 50 -257107
rect -50 -259325 50 -258325
rect -50 -260543 50 -259543
rect -50 -261761 50 -260761
rect -50 -262979 50 -261979
rect -50 -264197 50 -263197
rect -50 -265415 50 -264415
rect -50 -266633 50 -265633
rect -50 -267851 50 -266851
rect -50 -269069 50 -268069
rect -50 -270287 50 -269287
rect -50 -271505 50 -270505
rect -50 -272723 50 -271723
rect -50 -273941 50 -272941
rect -50 -275159 50 -274159
rect -50 -276377 50 -275377
rect -50 -277595 50 -276595
rect -50 -278813 50 -277813
rect -50 -280031 50 -279031
rect -50 -281249 50 -280249
rect -50 -282467 50 -281467
rect -50 -283685 50 -282685
rect -50 -284903 50 -283903
rect -50 -286121 50 -285121
rect -50 -287339 50 -286339
rect -50 -288557 50 -287557
rect -50 -289775 50 -288775
rect -50 -290993 50 -289993
rect -50 -292211 50 -291211
rect -50 -293429 50 -292429
rect -50 -294647 50 -293647
rect -50 -295865 50 -294865
rect -50 -297083 50 -296083
rect -50 -298301 50 -297301
rect -50 -299519 50 -298519
rect -50 -300737 50 -299737
rect -50 -301955 50 -300955
rect -50 -303173 50 -302173
rect -50 -304391 50 -303391
rect -50 -305609 50 -304609
rect -50 -306827 50 -305827
rect -50 -308045 50 -307045
rect -50 -309263 50 -308263
rect -50 -310481 50 -309481
rect -50 -311699 50 -310699
rect -50 -312917 50 -311917
rect -50 -314135 50 -313135
rect -50 -315353 50 -314353
rect -50 -316571 50 -315571
rect -50 -317789 50 -316789
rect -50 -319007 50 -318007
rect -50 -320225 50 -319225
rect -50 -321443 50 -320443
rect -50 -322661 50 -321661
rect -50 -323879 50 -322879
rect -50 -325097 50 -324097
rect -50 -326315 50 -325315
rect -50 -327533 50 -326533
rect -50 -328751 50 -327751
rect -50 -329969 50 -328969
rect -50 -331187 50 -330187
rect -50 -332405 50 -331405
rect -50 -333623 50 -332623
rect -50 -334841 50 -333841
rect -50 -336059 50 -335059
rect -50 -337277 50 -336277
rect -50 -338495 50 -337495
rect -50 -339713 50 -338713
rect -50 -340931 50 -339931
rect -50 -342149 50 -341149
rect -50 -343367 50 -342367
rect -50 -344585 50 -343585
rect -50 -345803 50 -344803
rect -50 -347021 50 -346021
rect -50 -348239 50 -347239
rect -50 -349457 50 -348457
rect -50 -350675 50 -349675
rect -50 -351893 50 -350893
rect -50 -353111 50 -352111
rect -50 -354329 50 -353329
rect -50 -355547 50 -354547
rect -50 -356765 50 -355765
rect -50 -357983 50 -356983
rect -50 -359201 50 -358201
rect -50 -360419 50 -359419
rect -50 -361637 50 -360637
rect -50 -362855 50 -361855
rect -50 -364073 50 -363073
rect -50 -365291 50 -364291
rect -50 -366509 50 -365509
rect -50 -367727 50 -366727
rect -50 -368945 50 -367945
rect -50 -370163 50 -369163
rect -50 -371381 50 -370381
rect -50 -372599 50 -371599
rect -50 -373817 50 -372817
rect -50 -375035 50 -374035
rect -50 -376253 50 -375253
rect -50 -377471 50 -376471
rect -50 -378689 50 -377689
rect -50 -379907 50 -378907
rect -50 -381125 50 -380125
rect -50 -382343 50 -381343
rect -50 -383561 50 -382561
rect -50 -384779 50 -383779
rect -50 -385997 50 -384997
rect -50 -387215 50 -386215
rect -50 -388433 50 -387433
rect -50 -389651 50 -388651
rect -50 -390869 50 -389869
rect -50 -392087 50 -391087
rect -50 -393305 50 -392305
rect -50 -394523 50 -393523
rect -50 -395741 50 -394741
rect -50 -396959 50 -395959
rect -50 -398177 50 -397177
rect -50 -399395 50 -398395
rect -50 -400613 50 -399613
rect -50 -401831 50 -400831
rect -50 -403049 50 -402049
rect -50 -404267 50 -403267
rect -50 -405485 50 -404485
rect -50 -406703 50 -405703
rect -50 -407921 50 -406921
rect -50 -409139 50 -408139
rect -50 -410357 50 -409357
rect -50 -411575 50 -410575
rect -50 -412793 50 -411793
rect -50 -414011 50 -413011
rect -50 -415229 50 -414229
rect -50 -416447 50 -415447
rect -50 -417665 50 -416665
rect -50 -418883 50 -417883
rect -50 -420101 50 -419101
rect -50 -421319 50 -420319
rect -50 -422537 50 -421537
rect -50 -423755 50 -422755
rect -50 -424973 50 -423973
rect -50 -426191 50 -425191
rect -50 -427409 50 -426409
rect -50 -428627 50 -427627
rect -50 -429845 50 -428845
rect -50 -431063 50 -430063
rect -50 -432281 50 -431281
rect -50 -433499 50 -432499
rect -50 -434717 50 -433717
rect -50 -435935 50 -434935
rect -50 -437153 50 -436153
rect -50 -438371 50 -437371
rect -50 -439589 50 -438589
rect -50 -440807 50 -439807
rect -50 -442025 50 -441025
rect -50 -443243 50 -442243
rect -50 -444461 50 -443461
rect -50 -445679 50 -444679
rect -50 -446897 50 -445897
rect -50 -448115 50 -447115
rect -50 -449333 50 -448333
rect -50 -450551 50 -449551
rect -50 -451769 50 -450769
rect -50 -452987 50 -451987
rect -50 -454205 50 -453205
rect -50 -455423 50 -454423
rect -50 -456641 50 -455641
rect -50 -457859 50 -456859
rect -50 -459077 50 -458077
rect -50 -460295 50 -459295
rect -50 -461513 50 -460513
rect -50 -462731 50 -461731
rect -50 -463949 50 -462949
rect -50 -465167 50 -464167
rect -50 -466385 50 -465385
rect -50 -467603 50 -466603
rect -50 -468821 50 -467821
rect -50 -470039 50 -469039
rect -50 -471257 50 -470257
rect -50 -472475 50 -471475
rect -50 -473693 50 -472693
rect -50 -474911 50 -473911
rect -50 -476129 50 -475129
rect -50 -477347 50 -476347
rect -50 -478565 50 -477565
rect -50 -479783 50 -478783
rect -50 -481001 50 -480001
rect -50 -482219 50 -481219
rect -50 -483437 50 -482437
rect -50 -484655 50 -483655
rect -50 -485873 50 -484873
rect -50 -487091 50 -486091
rect -50 -488309 50 -487309
rect -50 -489527 50 -488527
rect -50 -490745 50 -489745
rect -50 -491963 50 -490963
rect -50 -493181 50 -492181
rect -50 -494399 50 -493399
rect -50 -495617 50 -494617
rect -50 -496835 50 -495835
rect -50 -498053 50 -497053
rect -50 -499271 50 -498271
rect -50 -500489 50 -499489
rect -50 -501707 50 -500707
rect -50 -502925 50 -501925
rect -50 -504143 50 -503143
rect -50 -505361 50 -504361
rect -50 -506579 50 -505579
rect -50 -507797 50 -506797
rect -50 -509015 50 -508015
rect -50 -510233 50 -509233
rect -50 -511451 50 -510451
rect -50 -512669 50 -511669
rect -50 -513887 50 -512887
rect -50 -515105 50 -514105
rect -50 -516323 50 -515323
rect -50 -517541 50 -516541
rect -50 -518759 50 -517759
rect -50 -519977 50 -518977
rect -50 -521195 50 -520195
rect -50 -522413 50 -521413
rect -50 -523631 50 -522631
rect -50 -524849 50 -523849
rect -50 -526067 50 -525067
rect -50 -527285 50 -526285
rect -50 -528503 50 -527503
rect -50 -529721 50 -528721
rect -50 -530939 50 -529939
rect -50 -532157 50 -531157
rect -50 -533375 50 -532375
rect -50 -534593 50 -533593
rect -50 -535811 50 -534811
rect -50 -537029 50 -536029
rect -50 -538247 50 -537247
rect -50 -539465 50 -538465
rect -50 -540683 50 -539683
rect -50 -541901 50 -540901
rect -50 -543119 50 -542119
rect -50 -544337 50 -543337
rect -50 -545555 50 -544555
rect -50 -546773 50 -545773
rect -50 -547991 50 -546991
rect -50 -549209 50 -548209
rect -50 -550427 50 -549427
rect -50 -551645 50 -550645
rect -50 -552863 50 -551863
rect -50 -554081 50 -553081
rect -50 -555299 50 -554299
rect -50 -556517 50 -555517
rect -50 -557735 50 -556735
rect -50 -558953 50 -557953
rect -50 -560171 50 -559171
rect -50 -561389 50 -560389
rect -50 -562607 50 -561607
rect -50 -563825 50 -562825
rect -50 -565043 50 -564043
rect -50 -566261 50 -565261
rect -50 -567479 50 -566479
rect -50 -568697 50 -567697
rect -50 -569915 50 -568915
rect -50 -571133 50 -570133
rect -50 -572351 50 -571351
rect -50 -573569 50 -572569
rect -50 -574787 50 -573787
rect -50 -576005 50 -575005
rect -50 -577223 50 -576223
rect -50 -578441 50 -577441
rect -50 -579659 50 -578659
rect -50 -580877 50 -579877
rect -50 -582095 50 -581095
rect -50 -583313 50 -582313
rect -50 -584531 50 -583531
rect -50 -585749 50 -584749
rect -50 -586967 50 -585967
rect -50 -588185 50 -587185
rect -50 -589403 50 -588403
rect -50 -590621 50 -589621
rect -50 -591839 50 -590839
rect -50 -593057 50 -592057
rect -50 -594275 50 -593275
rect -50 -595493 50 -594493
rect -50 -596711 50 -595711
rect -50 -597929 50 -596929
rect -50 -599147 50 -598147
rect -50 -600365 50 -599365
rect -50 -601583 50 -600583
rect -50 -602801 50 -601801
rect -50 -604019 50 -603019
rect -50 -605237 50 -604237
rect -50 -606455 50 -605455
rect -50 -607673 50 -606673
rect -50 -608891 50 -607891
<< mvndiff >>
rect -108 608879 -50 608891
rect -108 607903 -96 608879
rect -62 607903 -50 608879
rect -108 607891 -50 607903
rect 50 608879 108 608891
rect 50 607903 62 608879
rect 96 607903 108 608879
rect 50 607891 108 607903
rect -108 607661 -50 607673
rect -108 606685 -96 607661
rect -62 606685 -50 607661
rect -108 606673 -50 606685
rect 50 607661 108 607673
rect 50 606685 62 607661
rect 96 606685 108 607661
rect 50 606673 108 606685
rect -108 606443 -50 606455
rect -108 605467 -96 606443
rect -62 605467 -50 606443
rect -108 605455 -50 605467
rect 50 606443 108 606455
rect 50 605467 62 606443
rect 96 605467 108 606443
rect 50 605455 108 605467
rect -108 605225 -50 605237
rect -108 604249 -96 605225
rect -62 604249 -50 605225
rect -108 604237 -50 604249
rect 50 605225 108 605237
rect 50 604249 62 605225
rect 96 604249 108 605225
rect 50 604237 108 604249
rect -108 604007 -50 604019
rect -108 603031 -96 604007
rect -62 603031 -50 604007
rect -108 603019 -50 603031
rect 50 604007 108 604019
rect 50 603031 62 604007
rect 96 603031 108 604007
rect 50 603019 108 603031
rect -108 602789 -50 602801
rect -108 601813 -96 602789
rect -62 601813 -50 602789
rect -108 601801 -50 601813
rect 50 602789 108 602801
rect 50 601813 62 602789
rect 96 601813 108 602789
rect 50 601801 108 601813
rect -108 601571 -50 601583
rect -108 600595 -96 601571
rect -62 600595 -50 601571
rect -108 600583 -50 600595
rect 50 601571 108 601583
rect 50 600595 62 601571
rect 96 600595 108 601571
rect 50 600583 108 600595
rect -108 600353 -50 600365
rect -108 599377 -96 600353
rect -62 599377 -50 600353
rect -108 599365 -50 599377
rect 50 600353 108 600365
rect 50 599377 62 600353
rect 96 599377 108 600353
rect 50 599365 108 599377
rect -108 599135 -50 599147
rect -108 598159 -96 599135
rect -62 598159 -50 599135
rect -108 598147 -50 598159
rect 50 599135 108 599147
rect 50 598159 62 599135
rect 96 598159 108 599135
rect 50 598147 108 598159
rect -108 597917 -50 597929
rect -108 596941 -96 597917
rect -62 596941 -50 597917
rect -108 596929 -50 596941
rect 50 597917 108 597929
rect 50 596941 62 597917
rect 96 596941 108 597917
rect 50 596929 108 596941
rect -108 596699 -50 596711
rect -108 595723 -96 596699
rect -62 595723 -50 596699
rect -108 595711 -50 595723
rect 50 596699 108 596711
rect 50 595723 62 596699
rect 96 595723 108 596699
rect 50 595711 108 595723
rect -108 595481 -50 595493
rect -108 594505 -96 595481
rect -62 594505 -50 595481
rect -108 594493 -50 594505
rect 50 595481 108 595493
rect 50 594505 62 595481
rect 96 594505 108 595481
rect 50 594493 108 594505
rect -108 594263 -50 594275
rect -108 593287 -96 594263
rect -62 593287 -50 594263
rect -108 593275 -50 593287
rect 50 594263 108 594275
rect 50 593287 62 594263
rect 96 593287 108 594263
rect 50 593275 108 593287
rect -108 593045 -50 593057
rect -108 592069 -96 593045
rect -62 592069 -50 593045
rect -108 592057 -50 592069
rect 50 593045 108 593057
rect 50 592069 62 593045
rect 96 592069 108 593045
rect 50 592057 108 592069
rect -108 591827 -50 591839
rect -108 590851 -96 591827
rect -62 590851 -50 591827
rect -108 590839 -50 590851
rect 50 591827 108 591839
rect 50 590851 62 591827
rect 96 590851 108 591827
rect 50 590839 108 590851
rect -108 590609 -50 590621
rect -108 589633 -96 590609
rect -62 589633 -50 590609
rect -108 589621 -50 589633
rect 50 590609 108 590621
rect 50 589633 62 590609
rect 96 589633 108 590609
rect 50 589621 108 589633
rect -108 589391 -50 589403
rect -108 588415 -96 589391
rect -62 588415 -50 589391
rect -108 588403 -50 588415
rect 50 589391 108 589403
rect 50 588415 62 589391
rect 96 588415 108 589391
rect 50 588403 108 588415
rect -108 588173 -50 588185
rect -108 587197 -96 588173
rect -62 587197 -50 588173
rect -108 587185 -50 587197
rect 50 588173 108 588185
rect 50 587197 62 588173
rect 96 587197 108 588173
rect 50 587185 108 587197
rect -108 586955 -50 586967
rect -108 585979 -96 586955
rect -62 585979 -50 586955
rect -108 585967 -50 585979
rect 50 586955 108 586967
rect 50 585979 62 586955
rect 96 585979 108 586955
rect 50 585967 108 585979
rect -108 585737 -50 585749
rect -108 584761 -96 585737
rect -62 584761 -50 585737
rect -108 584749 -50 584761
rect 50 585737 108 585749
rect 50 584761 62 585737
rect 96 584761 108 585737
rect 50 584749 108 584761
rect -108 584519 -50 584531
rect -108 583543 -96 584519
rect -62 583543 -50 584519
rect -108 583531 -50 583543
rect 50 584519 108 584531
rect 50 583543 62 584519
rect 96 583543 108 584519
rect 50 583531 108 583543
rect -108 583301 -50 583313
rect -108 582325 -96 583301
rect -62 582325 -50 583301
rect -108 582313 -50 582325
rect 50 583301 108 583313
rect 50 582325 62 583301
rect 96 582325 108 583301
rect 50 582313 108 582325
rect -108 582083 -50 582095
rect -108 581107 -96 582083
rect -62 581107 -50 582083
rect -108 581095 -50 581107
rect 50 582083 108 582095
rect 50 581107 62 582083
rect 96 581107 108 582083
rect 50 581095 108 581107
rect -108 580865 -50 580877
rect -108 579889 -96 580865
rect -62 579889 -50 580865
rect -108 579877 -50 579889
rect 50 580865 108 580877
rect 50 579889 62 580865
rect 96 579889 108 580865
rect 50 579877 108 579889
rect -108 579647 -50 579659
rect -108 578671 -96 579647
rect -62 578671 -50 579647
rect -108 578659 -50 578671
rect 50 579647 108 579659
rect 50 578671 62 579647
rect 96 578671 108 579647
rect 50 578659 108 578671
rect -108 578429 -50 578441
rect -108 577453 -96 578429
rect -62 577453 -50 578429
rect -108 577441 -50 577453
rect 50 578429 108 578441
rect 50 577453 62 578429
rect 96 577453 108 578429
rect 50 577441 108 577453
rect -108 577211 -50 577223
rect -108 576235 -96 577211
rect -62 576235 -50 577211
rect -108 576223 -50 576235
rect 50 577211 108 577223
rect 50 576235 62 577211
rect 96 576235 108 577211
rect 50 576223 108 576235
rect -108 575993 -50 576005
rect -108 575017 -96 575993
rect -62 575017 -50 575993
rect -108 575005 -50 575017
rect 50 575993 108 576005
rect 50 575017 62 575993
rect 96 575017 108 575993
rect 50 575005 108 575017
rect -108 574775 -50 574787
rect -108 573799 -96 574775
rect -62 573799 -50 574775
rect -108 573787 -50 573799
rect 50 574775 108 574787
rect 50 573799 62 574775
rect 96 573799 108 574775
rect 50 573787 108 573799
rect -108 573557 -50 573569
rect -108 572581 -96 573557
rect -62 572581 -50 573557
rect -108 572569 -50 572581
rect 50 573557 108 573569
rect 50 572581 62 573557
rect 96 572581 108 573557
rect 50 572569 108 572581
rect -108 572339 -50 572351
rect -108 571363 -96 572339
rect -62 571363 -50 572339
rect -108 571351 -50 571363
rect 50 572339 108 572351
rect 50 571363 62 572339
rect 96 571363 108 572339
rect 50 571351 108 571363
rect -108 571121 -50 571133
rect -108 570145 -96 571121
rect -62 570145 -50 571121
rect -108 570133 -50 570145
rect 50 571121 108 571133
rect 50 570145 62 571121
rect 96 570145 108 571121
rect 50 570133 108 570145
rect -108 569903 -50 569915
rect -108 568927 -96 569903
rect -62 568927 -50 569903
rect -108 568915 -50 568927
rect 50 569903 108 569915
rect 50 568927 62 569903
rect 96 568927 108 569903
rect 50 568915 108 568927
rect -108 568685 -50 568697
rect -108 567709 -96 568685
rect -62 567709 -50 568685
rect -108 567697 -50 567709
rect 50 568685 108 568697
rect 50 567709 62 568685
rect 96 567709 108 568685
rect 50 567697 108 567709
rect -108 567467 -50 567479
rect -108 566491 -96 567467
rect -62 566491 -50 567467
rect -108 566479 -50 566491
rect 50 567467 108 567479
rect 50 566491 62 567467
rect 96 566491 108 567467
rect 50 566479 108 566491
rect -108 566249 -50 566261
rect -108 565273 -96 566249
rect -62 565273 -50 566249
rect -108 565261 -50 565273
rect 50 566249 108 566261
rect 50 565273 62 566249
rect 96 565273 108 566249
rect 50 565261 108 565273
rect -108 565031 -50 565043
rect -108 564055 -96 565031
rect -62 564055 -50 565031
rect -108 564043 -50 564055
rect 50 565031 108 565043
rect 50 564055 62 565031
rect 96 564055 108 565031
rect 50 564043 108 564055
rect -108 563813 -50 563825
rect -108 562837 -96 563813
rect -62 562837 -50 563813
rect -108 562825 -50 562837
rect 50 563813 108 563825
rect 50 562837 62 563813
rect 96 562837 108 563813
rect 50 562825 108 562837
rect -108 562595 -50 562607
rect -108 561619 -96 562595
rect -62 561619 -50 562595
rect -108 561607 -50 561619
rect 50 562595 108 562607
rect 50 561619 62 562595
rect 96 561619 108 562595
rect 50 561607 108 561619
rect -108 561377 -50 561389
rect -108 560401 -96 561377
rect -62 560401 -50 561377
rect -108 560389 -50 560401
rect 50 561377 108 561389
rect 50 560401 62 561377
rect 96 560401 108 561377
rect 50 560389 108 560401
rect -108 560159 -50 560171
rect -108 559183 -96 560159
rect -62 559183 -50 560159
rect -108 559171 -50 559183
rect 50 560159 108 560171
rect 50 559183 62 560159
rect 96 559183 108 560159
rect 50 559171 108 559183
rect -108 558941 -50 558953
rect -108 557965 -96 558941
rect -62 557965 -50 558941
rect -108 557953 -50 557965
rect 50 558941 108 558953
rect 50 557965 62 558941
rect 96 557965 108 558941
rect 50 557953 108 557965
rect -108 557723 -50 557735
rect -108 556747 -96 557723
rect -62 556747 -50 557723
rect -108 556735 -50 556747
rect 50 557723 108 557735
rect 50 556747 62 557723
rect 96 556747 108 557723
rect 50 556735 108 556747
rect -108 556505 -50 556517
rect -108 555529 -96 556505
rect -62 555529 -50 556505
rect -108 555517 -50 555529
rect 50 556505 108 556517
rect 50 555529 62 556505
rect 96 555529 108 556505
rect 50 555517 108 555529
rect -108 555287 -50 555299
rect -108 554311 -96 555287
rect -62 554311 -50 555287
rect -108 554299 -50 554311
rect 50 555287 108 555299
rect 50 554311 62 555287
rect 96 554311 108 555287
rect 50 554299 108 554311
rect -108 554069 -50 554081
rect -108 553093 -96 554069
rect -62 553093 -50 554069
rect -108 553081 -50 553093
rect 50 554069 108 554081
rect 50 553093 62 554069
rect 96 553093 108 554069
rect 50 553081 108 553093
rect -108 552851 -50 552863
rect -108 551875 -96 552851
rect -62 551875 -50 552851
rect -108 551863 -50 551875
rect 50 552851 108 552863
rect 50 551875 62 552851
rect 96 551875 108 552851
rect 50 551863 108 551875
rect -108 551633 -50 551645
rect -108 550657 -96 551633
rect -62 550657 -50 551633
rect -108 550645 -50 550657
rect 50 551633 108 551645
rect 50 550657 62 551633
rect 96 550657 108 551633
rect 50 550645 108 550657
rect -108 550415 -50 550427
rect -108 549439 -96 550415
rect -62 549439 -50 550415
rect -108 549427 -50 549439
rect 50 550415 108 550427
rect 50 549439 62 550415
rect 96 549439 108 550415
rect 50 549427 108 549439
rect -108 549197 -50 549209
rect -108 548221 -96 549197
rect -62 548221 -50 549197
rect -108 548209 -50 548221
rect 50 549197 108 549209
rect 50 548221 62 549197
rect 96 548221 108 549197
rect 50 548209 108 548221
rect -108 547979 -50 547991
rect -108 547003 -96 547979
rect -62 547003 -50 547979
rect -108 546991 -50 547003
rect 50 547979 108 547991
rect 50 547003 62 547979
rect 96 547003 108 547979
rect 50 546991 108 547003
rect -108 546761 -50 546773
rect -108 545785 -96 546761
rect -62 545785 -50 546761
rect -108 545773 -50 545785
rect 50 546761 108 546773
rect 50 545785 62 546761
rect 96 545785 108 546761
rect 50 545773 108 545785
rect -108 545543 -50 545555
rect -108 544567 -96 545543
rect -62 544567 -50 545543
rect -108 544555 -50 544567
rect 50 545543 108 545555
rect 50 544567 62 545543
rect 96 544567 108 545543
rect 50 544555 108 544567
rect -108 544325 -50 544337
rect -108 543349 -96 544325
rect -62 543349 -50 544325
rect -108 543337 -50 543349
rect 50 544325 108 544337
rect 50 543349 62 544325
rect 96 543349 108 544325
rect 50 543337 108 543349
rect -108 543107 -50 543119
rect -108 542131 -96 543107
rect -62 542131 -50 543107
rect -108 542119 -50 542131
rect 50 543107 108 543119
rect 50 542131 62 543107
rect 96 542131 108 543107
rect 50 542119 108 542131
rect -108 541889 -50 541901
rect -108 540913 -96 541889
rect -62 540913 -50 541889
rect -108 540901 -50 540913
rect 50 541889 108 541901
rect 50 540913 62 541889
rect 96 540913 108 541889
rect 50 540901 108 540913
rect -108 540671 -50 540683
rect -108 539695 -96 540671
rect -62 539695 -50 540671
rect -108 539683 -50 539695
rect 50 540671 108 540683
rect 50 539695 62 540671
rect 96 539695 108 540671
rect 50 539683 108 539695
rect -108 539453 -50 539465
rect -108 538477 -96 539453
rect -62 538477 -50 539453
rect -108 538465 -50 538477
rect 50 539453 108 539465
rect 50 538477 62 539453
rect 96 538477 108 539453
rect 50 538465 108 538477
rect -108 538235 -50 538247
rect -108 537259 -96 538235
rect -62 537259 -50 538235
rect -108 537247 -50 537259
rect 50 538235 108 538247
rect 50 537259 62 538235
rect 96 537259 108 538235
rect 50 537247 108 537259
rect -108 537017 -50 537029
rect -108 536041 -96 537017
rect -62 536041 -50 537017
rect -108 536029 -50 536041
rect 50 537017 108 537029
rect 50 536041 62 537017
rect 96 536041 108 537017
rect 50 536029 108 536041
rect -108 535799 -50 535811
rect -108 534823 -96 535799
rect -62 534823 -50 535799
rect -108 534811 -50 534823
rect 50 535799 108 535811
rect 50 534823 62 535799
rect 96 534823 108 535799
rect 50 534811 108 534823
rect -108 534581 -50 534593
rect -108 533605 -96 534581
rect -62 533605 -50 534581
rect -108 533593 -50 533605
rect 50 534581 108 534593
rect 50 533605 62 534581
rect 96 533605 108 534581
rect 50 533593 108 533605
rect -108 533363 -50 533375
rect -108 532387 -96 533363
rect -62 532387 -50 533363
rect -108 532375 -50 532387
rect 50 533363 108 533375
rect 50 532387 62 533363
rect 96 532387 108 533363
rect 50 532375 108 532387
rect -108 532145 -50 532157
rect -108 531169 -96 532145
rect -62 531169 -50 532145
rect -108 531157 -50 531169
rect 50 532145 108 532157
rect 50 531169 62 532145
rect 96 531169 108 532145
rect 50 531157 108 531169
rect -108 530927 -50 530939
rect -108 529951 -96 530927
rect -62 529951 -50 530927
rect -108 529939 -50 529951
rect 50 530927 108 530939
rect 50 529951 62 530927
rect 96 529951 108 530927
rect 50 529939 108 529951
rect -108 529709 -50 529721
rect -108 528733 -96 529709
rect -62 528733 -50 529709
rect -108 528721 -50 528733
rect 50 529709 108 529721
rect 50 528733 62 529709
rect 96 528733 108 529709
rect 50 528721 108 528733
rect -108 528491 -50 528503
rect -108 527515 -96 528491
rect -62 527515 -50 528491
rect -108 527503 -50 527515
rect 50 528491 108 528503
rect 50 527515 62 528491
rect 96 527515 108 528491
rect 50 527503 108 527515
rect -108 527273 -50 527285
rect -108 526297 -96 527273
rect -62 526297 -50 527273
rect -108 526285 -50 526297
rect 50 527273 108 527285
rect 50 526297 62 527273
rect 96 526297 108 527273
rect 50 526285 108 526297
rect -108 526055 -50 526067
rect -108 525079 -96 526055
rect -62 525079 -50 526055
rect -108 525067 -50 525079
rect 50 526055 108 526067
rect 50 525079 62 526055
rect 96 525079 108 526055
rect 50 525067 108 525079
rect -108 524837 -50 524849
rect -108 523861 -96 524837
rect -62 523861 -50 524837
rect -108 523849 -50 523861
rect 50 524837 108 524849
rect 50 523861 62 524837
rect 96 523861 108 524837
rect 50 523849 108 523861
rect -108 523619 -50 523631
rect -108 522643 -96 523619
rect -62 522643 -50 523619
rect -108 522631 -50 522643
rect 50 523619 108 523631
rect 50 522643 62 523619
rect 96 522643 108 523619
rect 50 522631 108 522643
rect -108 522401 -50 522413
rect -108 521425 -96 522401
rect -62 521425 -50 522401
rect -108 521413 -50 521425
rect 50 522401 108 522413
rect 50 521425 62 522401
rect 96 521425 108 522401
rect 50 521413 108 521425
rect -108 521183 -50 521195
rect -108 520207 -96 521183
rect -62 520207 -50 521183
rect -108 520195 -50 520207
rect 50 521183 108 521195
rect 50 520207 62 521183
rect 96 520207 108 521183
rect 50 520195 108 520207
rect -108 519965 -50 519977
rect -108 518989 -96 519965
rect -62 518989 -50 519965
rect -108 518977 -50 518989
rect 50 519965 108 519977
rect 50 518989 62 519965
rect 96 518989 108 519965
rect 50 518977 108 518989
rect -108 518747 -50 518759
rect -108 517771 -96 518747
rect -62 517771 -50 518747
rect -108 517759 -50 517771
rect 50 518747 108 518759
rect 50 517771 62 518747
rect 96 517771 108 518747
rect 50 517759 108 517771
rect -108 517529 -50 517541
rect -108 516553 -96 517529
rect -62 516553 -50 517529
rect -108 516541 -50 516553
rect 50 517529 108 517541
rect 50 516553 62 517529
rect 96 516553 108 517529
rect 50 516541 108 516553
rect -108 516311 -50 516323
rect -108 515335 -96 516311
rect -62 515335 -50 516311
rect -108 515323 -50 515335
rect 50 516311 108 516323
rect 50 515335 62 516311
rect 96 515335 108 516311
rect 50 515323 108 515335
rect -108 515093 -50 515105
rect -108 514117 -96 515093
rect -62 514117 -50 515093
rect -108 514105 -50 514117
rect 50 515093 108 515105
rect 50 514117 62 515093
rect 96 514117 108 515093
rect 50 514105 108 514117
rect -108 513875 -50 513887
rect -108 512899 -96 513875
rect -62 512899 -50 513875
rect -108 512887 -50 512899
rect 50 513875 108 513887
rect 50 512899 62 513875
rect 96 512899 108 513875
rect 50 512887 108 512899
rect -108 512657 -50 512669
rect -108 511681 -96 512657
rect -62 511681 -50 512657
rect -108 511669 -50 511681
rect 50 512657 108 512669
rect 50 511681 62 512657
rect 96 511681 108 512657
rect 50 511669 108 511681
rect -108 511439 -50 511451
rect -108 510463 -96 511439
rect -62 510463 -50 511439
rect -108 510451 -50 510463
rect 50 511439 108 511451
rect 50 510463 62 511439
rect 96 510463 108 511439
rect 50 510451 108 510463
rect -108 510221 -50 510233
rect -108 509245 -96 510221
rect -62 509245 -50 510221
rect -108 509233 -50 509245
rect 50 510221 108 510233
rect 50 509245 62 510221
rect 96 509245 108 510221
rect 50 509233 108 509245
rect -108 509003 -50 509015
rect -108 508027 -96 509003
rect -62 508027 -50 509003
rect -108 508015 -50 508027
rect 50 509003 108 509015
rect 50 508027 62 509003
rect 96 508027 108 509003
rect 50 508015 108 508027
rect -108 507785 -50 507797
rect -108 506809 -96 507785
rect -62 506809 -50 507785
rect -108 506797 -50 506809
rect 50 507785 108 507797
rect 50 506809 62 507785
rect 96 506809 108 507785
rect 50 506797 108 506809
rect -108 506567 -50 506579
rect -108 505591 -96 506567
rect -62 505591 -50 506567
rect -108 505579 -50 505591
rect 50 506567 108 506579
rect 50 505591 62 506567
rect 96 505591 108 506567
rect 50 505579 108 505591
rect -108 505349 -50 505361
rect -108 504373 -96 505349
rect -62 504373 -50 505349
rect -108 504361 -50 504373
rect 50 505349 108 505361
rect 50 504373 62 505349
rect 96 504373 108 505349
rect 50 504361 108 504373
rect -108 504131 -50 504143
rect -108 503155 -96 504131
rect -62 503155 -50 504131
rect -108 503143 -50 503155
rect 50 504131 108 504143
rect 50 503155 62 504131
rect 96 503155 108 504131
rect 50 503143 108 503155
rect -108 502913 -50 502925
rect -108 501937 -96 502913
rect -62 501937 -50 502913
rect -108 501925 -50 501937
rect 50 502913 108 502925
rect 50 501937 62 502913
rect 96 501937 108 502913
rect 50 501925 108 501937
rect -108 501695 -50 501707
rect -108 500719 -96 501695
rect -62 500719 -50 501695
rect -108 500707 -50 500719
rect 50 501695 108 501707
rect 50 500719 62 501695
rect 96 500719 108 501695
rect 50 500707 108 500719
rect -108 500477 -50 500489
rect -108 499501 -96 500477
rect -62 499501 -50 500477
rect -108 499489 -50 499501
rect 50 500477 108 500489
rect 50 499501 62 500477
rect 96 499501 108 500477
rect 50 499489 108 499501
rect -108 499259 -50 499271
rect -108 498283 -96 499259
rect -62 498283 -50 499259
rect -108 498271 -50 498283
rect 50 499259 108 499271
rect 50 498283 62 499259
rect 96 498283 108 499259
rect 50 498271 108 498283
rect -108 498041 -50 498053
rect -108 497065 -96 498041
rect -62 497065 -50 498041
rect -108 497053 -50 497065
rect 50 498041 108 498053
rect 50 497065 62 498041
rect 96 497065 108 498041
rect 50 497053 108 497065
rect -108 496823 -50 496835
rect -108 495847 -96 496823
rect -62 495847 -50 496823
rect -108 495835 -50 495847
rect 50 496823 108 496835
rect 50 495847 62 496823
rect 96 495847 108 496823
rect 50 495835 108 495847
rect -108 495605 -50 495617
rect -108 494629 -96 495605
rect -62 494629 -50 495605
rect -108 494617 -50 494629
rect 50 495605 108 495617
rect 50 494629 62 495605
rect 96 494629 108 495605
rect 50 494617 108 494629
rect -108 494387 -50 494399
rect -108 493411 -96 494387
rect -62 493411 -50 494387
rect -108 493399 -50 493411
rect 50 494387 108 494399
rect 50 493411 62 494387
rect 96 493411 108 494387
rect 50 493399 108 493411
rect -108 493169 -50 493181
rect -108 492193 -96 493169
rect -62 492193 -50 493169
rect -108 492181 -50 492193
rect 50 493169 108 493181
rect 50 492193 62 493169
rect 96 492193 108 493169
rect 50 492181 108 492193
rect -108 491951 -50 491963
rect -108 490975 -96 491951
rect -62 490975 -50 491951
rect -108 490963 -50 490975
rect 50 491951 108 491963
rect 50 490975 62 491951
rect 96 490975 108 491951
rect 50 490963 108 490975
rect -108 490733 -50 490745
rect -108 489757 -96 490733
rect -62 489757 -50 490733
rect -108 489745 -50 489757
rect 50 490733 108 490745
rect 50 489757 62 490733
rect 96 489757 108 490733
rect 50 489745 108 489757
rect -108 489515 -50 489527
rect -108 488539 -96 489515
rect -62 488539 -50 489515
rect -108 488527 -50 488539
rect 50 489515 108 489527
rect 50 488539 62 489515
rect 96 488539 108 489515
rect 50 488527 108 488539
rect -108 488297 -50 488309
rect -108 487321 -96 488297
rect -62 487321 -50 488297
rect -108 487309 -50 487321
rect 50 488297 108 488309
rect 50 487321 62 488297
rect 96 487321 108 488297
rect 50 487309 108 487321
rect -108 487079 -50 487091
rect -108 486103 -96 487079
rect -62 486103 -50 487079
rect -108 486091 -50 486103
rect 50 487079 108 487091
rect 50 486103 62 487079
rect 96 486103 108 487079
rect 50 486091 108 486103
rect -108 485861 -50 485873
rect -108 484885 -96 485861
rect -62 484885 -50 485861
rect -108 484873 -50 484885
rect 50 485861 108 485873
rect 50 484885 62 485861
rect 96 484885 108 485861
rect 50 484873 108 484885
rect -108 484643 -50 484655
rect -108 483667 -96 484643
rect -62 483667 -50 484643
rect -108 483655 -50 483667
rect 50 484643 108 484655
rect 50 483667 62 484643
rect 96 483667 108 484643
rect 50 483655 108 483667
rect -108 483425 -50 483437
rect -108 482449 -96 483425
rect -62 482449 -50 483425
rect -108 482437 -50 482449
rect 50 483425 108 483437
rect 50 482449 62 483425
rect 96 482449 108 483425
rect 50 482437 108 482449
rect -108 482207 -50 482219
rect -108 481231 -96 482207
rect -62 481231 -50 482207
rect -108 481219 -50 481231
rect 50 482207 108 482219
rect 50 481231 62 482207
rect 96 481231 108 482207
rect 50 481219 108 481231
rect -108 480989 -50 481001
rect -108 480013 -96 480989
rect -62 480013 -50 480989
rect -108 480001 -50 480013
rect 50 480989 108 481001
rect 50 480013 62 480989
rect 96 480013 108 480989
rect 50 480001 108 480013
rect -108 479771 -50 479783
rect -108 478795 -96 479771
rect -62 478795 -50 479771
rect -108 478783 -50 478795
rect 50 479771 108 479783
rect 50 478795 62 479771
rect 96 478795 108 479771
rect 50 478783 108 478795
rect -108 478553 -50 478565
rect -108 477577 -96 478553
rect -62 477577 -50 478553
rect -108 477565 -50 477577
rect 50 478553 108 478565
rect 50 477577 62 478553
rect 96 477577 108 478553
rect 50 477565 108 477577
rect -108 477335 -50 477347
rect -108 476359 -96 477335
rect -62 476359 -50 477335
rect -108 476347 -50 476359
rect 50 477335 108 477347
rect 50 476359 62 477335
rect 96 476359 108 477335
rect 50 476347 108 476359
rect -108 476117 -50 476129
rect -108 475141 -96 476117
rect -62 475141 -50 476117
rect -108 475129 -50 475141
rect 50 476117 108 476129
rect 50 475141 62 476117
rect 96 475141 108 476117
rect 50 475129 108 475141
rect -108 474899 -50 474911
rect -108 473923 -96 474899
rect -62 473923 -50 474899
rect -108 473911 -50 473923
rect 50 474899 108 474911
rect 50 473923 62 474899
rect 96 473923 108 474899
rect 50 473911 108 473923
rect -108 473681 -50 473693
rect -108 472705 -96 473681
rect -62 472705 -50 473681
rect -108 472693 -50 472705
rect 50 473681 108 473693
rect 50 472705 62 473681
rect 96 472705 108 473681
rect 50 472693 108 472705
rect -108 472463 -50 472475
rect -108 471487 -96 472463
rect -62 471487 -50 472463
rect -108 471475 -50 471487
rect 50 472463 108 472475
rect 50 471487 62 472463
rect 96 471487 108 472463
rect 50 471475 108 471487
rect -108 471245 -50 471257
rect -108 470269 -96 471245
rect -62 470269 -50 471245
rect -108 470257 -50 470269
rect 50 471245 108 471257
rect 50 470269 62 471245
rect 96 470269 108 471245
rect 50 470257 108 470269
rect -108 470027 -50 470039
rect -108 469051 -96 470027
rect -62 469051 -50 470027
rect -108 469039 -50 469051
rect 50 470027 108 470039
rect 50 469051 62 470027
rect 96 469051 108 470027
rect 50 469039 108 469051
rect -108 468809 -50 468821
rect -108 467833 -96 468809
rect -62 467833 -50 468809
rect -108 467821 -50 467833
rect 50 468809 108 468821
rect 50 467833 62 468809
rect 96 467833 108 468809
rect 50 467821 108 467833
rect -108 467591 -50 467603
rect -108 466615 -96 467591
rect -62 466615 -50 467591
rect -108 466603 -50 466615
rect 50 467591 108 467603
rect 50 466615 62 467591
rect 96 466615 108 467591
rect 50 466603 108 466615
rect -108 466373 -50 466385
rect -108 465397 -96 466373
rect -62 465397 -50 466373
rect -108 465385 -50 465397
rect 50 466373 108 466385
rect 50 465397 62 466373
rect 96 465397 108 466373
rect 50 465385 108 465397
rect -108 465155 -50 465167
rect -108 464179 -96 465155
rect -62 464179 -50 465155
rect -108 464167 -50 464179
rect 50 465155 108 465167
rect 50 464179 62 465155
rect 96 464179 108 465155
rect 50 464167 108 464179
rect -108 463937 -50 463949
rect -108 462961 -96 463937
rect -62 462961 -50 463937
rect -108 462949 -50 462961
rect 50 463937 108 463949
rect 50 462961 62 463937
rect 96 462961 108 463937
rect 50 462949 108 462961
rect -108 462719 -50 462731
rect -108 461743 -96 462719
rect -62 461743 -50 462719
rect -108 461731 -50 461743
rect 50 462719 108 462731
rect 50 461743 62 462719
rect 96 461743 108 462719
rect 50 461731 108 461743
rect -108 461501 -50 461513
rect -108 460525 -96 461501
rect -62 460525 -50 461501
rect -108 460513 -50 460525
rect 50 461501 108 461513
rect 50 460525 62 461501
rect 96 460525 108 461501
rect 50 460513 108 460525
rect -108 460283 -50 460295
rect -108 459307 -96 460283
rect -62 459307 -50 460283
rect -108 459295 -50 459307
rect 50 460283 108 460295
rect 50 459307 62 460283
rect 96 459307 108 460283
rect 50 459295 108 459307
rect -108 459065 -50 459077
rect -108 458089 -96 459065
rect -62 458089 -50 459065
rect -108 458077 -50 458089
rect 50 459065 108 459077
rect 50 458089 62 459065
rect 96 458089 108 459065
rect 50 458077 108 458089
rect -108 457847 -50 457859
rect -108 456871 -96 457847
rect -62 456871 -50 457847
rect -108 456859 -50 456871
rect 50 457847 108 457859
rect 50 456871 62 457847
rect 96 456871 108 457847
rect 50 456859 108 456871
rect -108 456629 -50 456641
rect -108 455653 -96 456629
rect -62 455653 -50 456629
rect -108 455641 -50 455653
rect 50 456629 108 456641
rect 50 455653 62 456629
rect 96 455653 108 456629
rect 50 455641 108 455653
rect -108 455411 -50 455423
rect -108 454435 -96 455411
rect -62 454435 -50 455411
rect -108 454423 -50 454435
rect 50 455411 108 455423
rect 50 454435 62 455411
rect 96 454435 108 455411
rect 50 454423 108 454435
rect -108 454193 -50 454205
rect -108 453217 -96 454193
rect -62 453217 -50 454193
rect -108 453205 -50 453217
rect 50 454193 108 454205
rect 50 453217 62 454193
rect 96 453217 108 454193
rect 50 453205 108 453217
rect -108 452975 -50 452987
rect -108 451999 -96 452975
rect -62 451999 -50 452975
rect -108 451987 -50 451999
rect 50 452975 108 452987
rect 50 451999 62 452975
rect 96 451999 108 452975
rect 50 451987 108 451999
rect -108 451757 -50 451769
rect -108 450781 -96 451757
rect -62 450781 -50 451757
rect -108 450769 -50 450781
rect 50 451757 108 451769
rect 50 450781 62 451757
rect 96 450781 108 451757
rect 50 450769 108 450781
rect -108 450539 -50 450551
rect -108 449563 -96 450539
rect -62 449563 -50 450539
rect -108 449551 -50 449563
rect 50 450539 108 450551
rect 50 449563 62 450539
rect 96 449563 108 450539
rect 50 449551 108 449563
rect -108 449321 -50 449333
rect -108 448345 -96 449321
rect -62 448345 -50 449321
rect -108 448333 -50 448345
rect 50 449321 108 449333
rect 50 448345 62 449321
rect 96 448345 108 449321
rect 50 448333 108 448345
rect -108 448103 -50 448115
rect -108 447127 -96 448103
rect -62 447127 -50 448103
rect -108 447115 -50 447127
rect 50 448103 108 448115
rect 50 447127 62 448103
rect 96 447127 108 448103
rect 50 447115 108 447127
rect -108 446885 -50 446897
rect -108 445909 -96 446885
rect -62 445909 -50 446885
rect -108 445897 -50 445909
rect 50 446885 108 446897
rect 50 445909 62 446885
rect 96 445909 108 446885
rect 50 445897 108 445909
rect -108 445667 -50 445679
rect -108 444691 -96 445667
rect -62 444691 -50 445667
rect -108 444679 -50 444691
rect 50 445667 108 445679
rect 50 444691 62 445667
rect 96 444691 108 445667
rect 50 444679 108 444691
rect -108 444449 -50 444461
rect -108 443473 -96 444449
rect -62 443473 -50 444449
rect -108 443461 -50 443473
rect 50 444449 108 444461
rect 50 443473 62 444449
rect 96 443473 108 444449
rect 50 443461 108 443473
rect -108 443231 -50 443243
rect -108 442255 -96 443231
rect -62 442255 -50 443231
rect -108 442243 -50 442255
rect 50 443231 108 443243
rect 50 442255 62 443231
rect 96 442255 108 443231
rect 50 442243 108 442255
rect -108 442013 -50 442025
rect -108 441037 -96 442013
rect -62 441037 -50 442013
rect -108 441025 -50 441037
rect 50 442013 108 442025
rect 50 441037 62 442013
rect 96 441037 108 442013
rect 50 441025 108 441037
rect -108 440795 -50 440807
rect -108 439819 -96 440795
rect -62 439819 -50 440795
rect -108 439807 -50 439819
rect 50 440795 108 440807
rect 50 439819 62 440795
rect 96 439819 108 440795
rect 50 439807 108 439819
rect -108 439577 -50 439589
rect -108 438601 -96 439577
rect -62 438601 -50 439577
rect -108 438589 -50 438601
rect 50 439577 108 439589
rect 50 438601 62 439577
rect 96 438601 108 439577
rect 50 438589 108 438601
rect -108 438359 -50 438371
rect -108 437383 -96 438359
rect -62 437383 -50 438359
rect -108 437371 -50 437383
rect 50 438359 108 438371
rect 50 437383 62 438359
rect 96 437383 108 438359
rect 50 437371 108 437383
rect -108 437141 -50 437153
rect -108 436165 -96 437141
rect -62 436165 -50 437141
rect -108 436153 -50 436165
rect 50 437141 108 437153
rect 50 436165 62 437141
rect 96 436165 108 437141
rect 50 436153 108 436165
rect -108 435923 -50 435935
rect -108 434947 -96 435923
rect -62 434947 -50 435923
rect -108 434935 -50 434947
rect 50 435923 108 435935
rect 50 434947 62 435923
rect 96 434947 108 435923
rect 50 434935 108 434947
rect -108 434705 -50 434717
rect -108 433729 -96 434705
rect -62 433729 -50 434705
rect -108 433717 -50 433729
rect 50 434705 108 434717
rect 50 433729 62 434705
rect 96 433729 108 434705
rect 50 433717 108 433729
rect -108 433487 -50 433499
rect -108 432511 -96 433487
rect -62 432511 -50 433487
rect -108 432499 -50 432511
rect 50 433487 108 433499
rect 50 432511 62 433487
rect 96 432511 108 433487
rect 50 432499 108 432511
rect -108 432269 -50 432281
rect -108 431293 -96 432269
rect -62 431293 -50 432269
rect -108 431281 -50 431293
rect 50 432269 108 432281
rect 50 431293 62 432269
rect 96 431293 108 432269
rect 50 431281 108 431293
rect -108 431051 -50 431063
rect -108 430075 -96 431051
rect -62 430075 -50 431051
rect -108 430063 -50 430075
rect 50 431051 108 431063
rect 50 430075 62 431051
rect 96 430075 108 431051
rect 50 430063 108 430075
rect -108 429833 -50 429845
rect -108 428857 -96 429833
rect -62 428857 -50 429833
rect -108 428845 -50 428857
rect 50 429833 108 429845
rect 50 428857 62 429833
rect 96 428857 108 429833
rect 50 428845 108 428857
rect -108 428615 -50 428627
rect -108 427639 -96 428615
rect -62 427639 -50 428615
rect -108 427627 -50 427639
rect 50 428615 108 428627
rect 50 427639 62 428615
rect 96 427639 108 428615
rect 50 427627 108 427639
rect -108 427397 -50 427409
rect -108 426421 -96 427397
rect -62 426421 -50 427397
rect -108 426409 -50 426421
rect 50 427397 108 427409
rect 50 426421 62 427397
rect 96 426421 108 427397
rect 50 426409 108 426421
rect -108 426179 -50 426191
rect -108 425203 -96 426179
rect -62 425203 -50 426179
rect -108 425191 -50 425203
rect 50 426179 108 426191
rect 50 425203 62 426179
rect 96 425203 108 426179
rect 50 425191 108 425203
rect -108 424961 -50 424973
rect -108 423985 -96 424961
rect -62 423985 -50 424961
rect -108 423973 -50 423985
rect 50 424961 108 424973
rect 50 423985 62 424961
rect 96 423985 108 424961
rect 50 423973 108 423985
rect -108 423743 -50 423755
rect -108 422767 -96 423743
rect -62 422767 -50 423743
rect -108 422755 -50 422767
rect 50 423743 108 423755
rect 50 422767 62 423743
rect 96 422767 108 423743
rect 50 422755 108 422767
rect -108 422525 -50 422537
rect -108 421549 -96 422525
rect -62 421549 -50 422525
rect -108 421537 -50 421549
rect 50 422525 108 422537
rect 50 421549 62 422525
rect 96 421549 108 422525
rect 50 421537 108 421549
rect -108 421307 -50 421319
rect -108 420331 -96 421307
rect -62 420331 -50 421307
rect -108 420319 -50 420331
rect 50 421307 108 421319
rect 50 420331 62 421307
rect 96 420331 108 421307
rect 50 420319 108 420331
rect -108 420089 -50 420101
rect -108 419113 -96 420089
rect -62 419113 -50 420089
rect -108 419101 -50 419113
rect 50 420089 108 420101
rect 50 419113 62 420089
rect 96 419113 108 420089
rect 50 419101 108 419113
rect -108 418871 -50 418883
rect -108 417895 -96 418871
rect -62 417895 -50 418871
rect -108 417883 -50 417895
rect 50 418871 108 418883
rect 50 417895 62 418871
rect 96 417895 108 418871
rect 50 417883 108 417895
rect -108 417653 -50 417665
rect -108 416677 -96 417653
rect -62 416677 -50 417653
rect -108 416665 -50 416677
rect 50 417653 108 417665
rect 50 416677 62 417653
rect 96 416677 108 417653
rect 50 416665 108 416677
rect -108 416435 -50 416447
rect -108 415459 -96 416435
rect -62 415459 -50 416435
rect -108 415447 -50 415459
rect 50 416435 108 416447
rect 50 415459 62 416435
rect 96 415459 108 416435
rect 50 415447 108 415459
rect -108 415217 -50 415229
rect -108 414241 -96 415217
rect -62 414241 -50 415217
rect -108 414229 -50 414241
rect 50 415217 108 415229
rect 50 414241 62 415217
rect 96 414241 108 415217
rect 50 414229 108 414241
rect -108 413999 -50 414011
rect -108 413023 -96 413999
rect -62 413023 -50 413999
rect -108 413011 -50 413023
rect 50 413999 108 414011
rect 50 413023 62 413999
rect 96 413023 108 413999
rect 50 413011 108 413023
rect -108 412781 -50 412793
rect -108 411805 -96 412781
rect -62 411805 -50 412781
rect -108 411793 -50 411805
rect 50 412781 108 412793
rect 50 411805 62 412781
rect 96 411805 108 412781
rect 50 411793 108 411805
rect -108 411563 -50 411575
rect -108 410587 -96 411563
rect -62 410587 -50 411563
rect -108 410575 -50 410587
rect 50 411563 108 411575
rect 50 410587 62 411563
rect 96 410587 108 411563
rect 50 410575 108 410587
rect -108 410345 -50 410357
rect -108 409369 -96 410345
rect -62 409369 -50 410345
rect -108 409357 -50 409369
rect 50 410345 108 410357
rect 50 409369 62 410345
rect 96 409369 108 410345
rect 50 409357 108 409369
rect -108 409127 -50 409139
rect -108 408151 -96 409127
rect -62 408151 -50 409127
rect -108 408139 -50 408151
rect 50 409127 108 409139
rect 50 408151 62 409127
rect 96 408151 108 409127
rect 50 408139 108 408151
rect -108 407909 -50 407921
rect -108 406933 -96 407909
rect -62 406933 -50 407909
rect -108 406921 -50 406933
rect 50 407909 108 407921
rect 50 406933 62 407909
rect 96 406933 108 407909
rect 50 406921 108 406933
rect -108 406691 -50 406703
rect -108 405715 -96 406691
rect -62 405715 -50 406691
rect -108 405703 -50 405715
rect 50 406691 108 406703
rect 50 405715 62 406691
rect 96 405715 108 406691
rect 50 405703 108 405715
rect -108 405473 -50 405485
rect -108 404497 -96 405473
rect -62 404497 -50 405473
rect -108 404485 -50 404497
rect 50 405473 108 405485
rect 50 404497 62 405473
rect 96 404497 108 405473
rect 50 404485 108 404497
rect -108 404255 -50 404267
rect -108 403279 -96 404255
rect -62 403279 -50 404255
rect -108 403267 -50 403279
rect 50 404255 108 404267
rect 50 403279 62 404255
rect 96 403279 108 404255
rect 50 403267 108 403279
rect -108 403037 -50 403049
rect -108 402061 -96 403037
rect -62 402061 -50 403037
rect -108 402049 -50 402061
rect 50 403037 108 403049
rect 50 402061 62 403037
rect 96 402061 108 403037
rect 50 402049 108 402061
rect -108 401819 -50 401831
rect -108 400843 -96 401819
rect -62 400843 -50 401819
rect -108 400831 -50 400843
rect 50 401819 108 401831
rect 50 400843 62 401819
rect 96 400843 108 401819
rect 50 400831 108 400843
rect -108 400601 -50 400613
rect -108 399625 -96 400601
rect -62 399625 -50 400601
rect -108 399613 -50 399625
rect 50 400601 108 400613
rect 50 399625 62 400601
rect 96 399625 108 400601
rect 50 399613 108 399625
rect -108 399383 -50 399395
rect -108 398407 -96 399383
rect -62 398407 -50 399383
rect -108 398395 -50 398407
rect 50 399383 108 399395
rect 50 398407 62 399383
rect 96 398407 108 399383
rect 50 398395 108 398407
rect -108 398165 -50 398177
rect -108 397189 -96 398165
rect -62 397189 -50 398165
rect -108 397177 -50 397189
rect 50 398165 108 398177
rect 50 397189 62 398165
rect 96 397189 108 398165
rect 50 397177 108 397189
rect -108 396947 -50 396959
rect -108 395971 -96 396947
rect -62 395971 -50 396947
rect -108 395959 -50 395971
rect 50 396947 108 396959
rect 50 395971 62 396947
rect 96 395971 108 396947
rect 50 395959 108 395971
rect -108 395729 -50 395741
rect -108 394753 -96 395729
rect -62 394753 -50 395729
rect -108 394741 -50 394753
rect 50 395729 108 395741
rect 50 394753 62 395729
rect 96 394753 108 395729
rect 50 394741 108 394753
rect -108 394511 -50 394523
rect -108 393535 -96 394511
rect -62 393535 -50 394511
rect -108 393523 -50 393535
rect 50 394511 108 394523
rect 50 393535 62 394511
rect 96 393535 108 394511
rect 50 393523 108 393535
rect -108 393293 -50 393305
rect -108 392317 -96 393293
rect -62 392317 -50 393293
rect -108 392305 -50 392317
rect 50 393293 108 393305
rect 50 392317 62 393293
rect 96 392317 108 393293
rect 50 392305 108 392317
rect -108 392075 -50 392087
rect -108 391099 -96 392075
rect -62 391099 -50 392075
rect -108 391087 -50 391099
rect 50 392075 108 392087
rect 50 391099 62 392075
rect 96 391099 108 392075
rect 50 391087 108 391099
rect -108 390857 -50 390869
rect -108 389881 -96 390857
rect -62 389881 -50 390857
rect -108 389869 -50 389881
rect 50 390857 108 390869
rect 50 389881 62 390857
rect 96 389881 108 390857
rect 50 389869 108 389881
rect -108 389639 -50 389651
rect -108 388663 -96 389639
rect -62 388663 -50 389639
rect -108 388651 -50 388663
rect 50 389639 108 389651
rect 50 388663 62 389639
rect 96 388663 108 389639
rect 50 388651 108 388663
rect -108 388421 -50 388433
rect -108 387445 -96 388421
rect -62 387445 -50 388421
rect -108 387433 -50 387445
rect 50 388421 108 388433
rect 50 387445 62 388421
rect 96 387445 108 388421
rect 50 387433 108 387445
rect -108 387203 -50 387215
rect -108 386227 -96 387203
rect -62 386227 -50 387203
rect -108 386215 -50 386227
rect 50 387203 108 387215
rect 50 386227 62 387203
rect 96 386227 108 387203
rect 50 386215 108 386227
rect -108 385985 -50 385997
rect -108 385009 -96 385985
rect -62 385009 -50 385985
rect -108 384997 -50 385009
rect 50 385985 108 385997
rect 50 385009 62 385985
rect 96 385009 108 385985
rect 50 384997 108 385009
rect -108 384767 -50 384779
rect -108 383791 -96 384767
rect -62 383791 -50 384767
rect -108 383779 -50 383791
rect 50 384767 108 384779
rect 50 383791 62 384767
rect 96 383791 108 384767
rect 50 383779 108 383791
rect -108 383549 -50 383561
rect -108 382573 -96 383549
rect -62 382573 -50 383549
rect -108 382561 -50 382573
rect 50 383549 108 383561
rect 50 382573 62 383549
rect 96 382573 108 383549
rect 50 382561 108 382573
rect -108 382331 -50 382343
rect -108 381355 -96 382331
rect -62 381355 -50 382331
rect -108 381343 -50 381355
rect 50 382331 108 382343
rect 50 381355 62 382331
rect 96 381355 108 382331
rect 50 381343 108 381355
rect -108 381113 -50 381125
rect -108 380137 -96 381113
rect -62 380137 -50 381113
rect -108 380125 -50 380137
rect 50 381113 108 381125
rect 50 380137 62 381113
rect 96 380137 108 381113
rect 50 380125 108 380137
rect -108 379895 -50 379907
rect -108 378919 -96 379895
rect -62 378919 -50 379895
rect -108 378907 -50 378919
rect 50 379895 108 379907
rect 50 378919 62 379895
rect 96 378919 108 379895
rect 50 378907 108 378919
rect -108 378677 -50 378689
rect -108 377701 -96 378677
rect -62 377701 -50 378677
rect -108 377689 -50 377701
rect 50 378677 108 378689
rect 50 377701 62 378677
rect 96 377701 108 378677
rect 50 377689 108 377701
rect -108 377459 -50 377471
rect -108 376483 -96 377459
rect -62 376483 -50 377459
rect -108 376471 -50 376483
rect 50 377459 108 377471
rect 50 376483 62 377459
rect 96 376483 108 377459
rect 50 376471 108 376483
rect -108 376241 -50 376253
rect -108 375265 -96 376241
rect -62 375265 -50 376241
rect -108 375253 -50 375265
rect 50 376241 108 376253
rect 50 375265 62 376241
rect 96 375265 108 376241
rect 50 375253 108 375265
rect -108 375023 -50 375035
rect -108 374047 -96 375023
rect -62 374047 -50 375023
rect -108 374035 -50 374047
rect 50 375023 108 375035
rect 50 374047 62 375023
rect 96 374047 108 375023
rect 50 374035 108 374047
rect -108 373805 -50 373817
rect -108 372829 -96 373805
rect -62 372829 -50 373805
rect -108 372817 -50 372829
rect 50 373805 108 373817
rect 50 372829 62 373805
rect 96 372829 108 373805
rect 50 372817 108 372829
rect -108 372587 -50 372599
rect -108 371611 -96 372587
rect -62 371611 -50 372587
rect -108 371599 -50 371611
rect 50 372587 108 372599
rect 50 371611 62 372587
rect 96 371611 108 372587
rect 50 371599 108 371611
rect -108 371369 -50 371381
rect -108 370393 -96 371369
rect -62 370393 -50 371369
rect -108 370381 -50 370393
rect 50 371369 108 371381
rect 50 370393 62 371369
rect 96 370393 108 371369
rect 50 370381 108 370393
rect -108 370151 -50 370163
rect -108 369175 -96 370151
rect -62 369175 -50 370151
rect -108 369163 -50 369175
rect 50 370151 108 370163
rect 50 369175 62 370151
rect 96 369175 108 370151
rect 50 369163 108 369175
rect -108 368933 -50 368945
rect -108 367957 -96 368933
rect -62 367957 -50 368933
rect -108 367945 -50 367957
rect 50 368933 108 368945
rect 50 367957 62 368933
rect 96 367957 108 368933
rect 50 367945 108 367957
rect -108 367715 -50 367727
rect -108 366739 -96 367715
rect -62 366739 -50 367715
rect -108 366727 -50 366739
rect 50 367715 108 367727
rect 50 366739 62 367715
rect 96 366739 108 367715
rect 50 366727 108 366739
rect -108 366497 -50 366509
rect -108 365521 -96 366497
rect -62 365521 -50 366497
rect -108 365509 -50 365521
rect 50 366497 108 366509
rect 50 365521 62 366497
rect 96 365521 108 366497
rect 50 365509 108 365521
rect -108 365279 -50 365291
rect -108 364303 -96 365279
rect -62 364303 -50 365279
rect -108 364291 -50 364303
rect 50 365279 108 365291
rect 50 364303 62 365279
rect 96 364303 108 365279
rect 50 364291 108 364303
rect -108 364061 -50 364073
rect -108 363085 -96 364061
rect -62 363085 -50 364061
rect -108 363073 -50 363085
rect 50 364061 108 364073
rect 50 363085 62 364061
rect 96 363085 108 364061
rect 50 363073 108 363085
rect -108 362843 -50 362855
rect -108 361867 -96 362843
rect -62 361867 -50 362843
rect -108 361855 -50 361867
rect 50 362843 108 362855
rect 50 361867 62 362843
rect 96 361867 108 362843
rect 50 361855 108 361867
rect -108 361625 -50 361637
rect -108 360649 -96 361625
rect -62 360649 -50 361625
rect -108 360637 -50 360649
rect 50 361625 108 361637
rect 50 360649 62 361625
rect 96 360649 108 361625
rect 50 360637 108 360649
rect -108 360407 -50 360419
rect -108 359431 -96 360407
rect -62 359431 -50 360407
rect -108 359419 -50 359431
rect 50 360407 108 360419
rect 50 359431 62 360407
rect 96 359431 108 360407
rect 50 359419 108 359431
rect -108 359189 -50 359201
rect -108 358213 -96 359189
rect -62 358213 -50 359189
rect -108 358201 -50 358213
rect 50 359189 108 359201
rect 50 358213 62 359189
rect 96 358213 108 359189
rect 50 358201 108 358213
rect -108 357971 -50 357983
rect -108 356995 -96 357971
rect -62 356995 -50 357971
rect -108 356983 -50 356995
rect 50 357971 108 357983
rect 50 356995 62 357971
rect 96 356995 108 357971
rect 50 356983 108 356995
rect -108 356753 -50 356765
rect -108 355777 -96 356753
rect -62 355777 -50 356753
rect -108 355765 -50 355777
rect 50 356753 108 356765
rect 50 355777 62 356753
rect 96 355777 108 356753
rect 50 355765 108 355777
rect -108 355535 -50 355547
rect -108 354559 -96 355535
rect -62 354559 -50 355535
rect -108 354547 -50 354559
rect 50 355535 108 355547
rect 50 354559 62 355535
rect 96 354559 108 355535
rect 50 354547 108 354559
rect -108 354317 -50 354329
rect -108 353341 -96 354317
rect -62 353341 -50 354317
rect -108 353329 -50 353341
rect 50 354317 108 354329
rect 50 353341 62 354317
rect 96 353341 108 354317
rect 50 353329 108 353341
rect -108 353099 -50 353111
rect -108 352123 -96 353099
rect -62 352123 -50 353099
rect -108 352111 -50 352123
rect 50 353099 108 353111
rect 50 352123 62 353099
rect 96 352123 108 353099
rect 50 352111 108 352123
rect -108 351881 -50 351893
rect -108 350905 -96 351881
rect -62 350905 -50 351881
rect -108 350893 -50 350905
rect 50 351881 108 351893
rect 50 350905 62 351881
rect 96 350905 108 351881
rect 50 350893 108 350905
rect -108 350663 -50 350675
rect -108 349687 -96 350663
rect -62 349687 -50 350663
rect -108 349675 -50 349687
rect 50 350663 108 350675
rect 50 349687 62 350663
rect 96 349687 108 350663
rect 50 349675 108 349687
rect -108 349445 -50 349457
rect -108 348469 -96 349445
rect -62 348469 -50 349445
rect -108 348457 -50 348469
rect 50 349445 108 349457
rect 50 348469 62 349445
rect 96 348469 108 349445
rect 50 348457 108 348469
rect -108 348227 -50 348239
rect -108 347251 -96 348227
rect -62 347251 -50 348227
rect -108 347239 -50 347251
rect 50 348227 108 348239
rect 50 347251 62 348227
rect 96 347251 108 348227
rect 50 347239 108 347251
rect -108 347009 -50 347021
rect -108 346033 -96 347009
rect -62 346033 -50 347009
rect -108 346021 -50 346033
rect 50 347009 108 347021
rect 50 346033 62 347009
rect 96 346033 108 347009
rect 50 346021 108 346033
rect -108 345791 -50 345803
rect -108 344815 -96 345791
rect -62 344815 -50 345791
rect -108 344803 -50 344815
rect 50 345791 108 345803
rect 50 344815 62 345791
rect 96 344815 108 345791
rect 50 344803 108 344815
rect -108 344573 -50 344585
rect -108 343597 -96 344573
rect -62 343597 -50 344573
rect -108 343585 -50 343597
rect 50 344573 108 344585
rect 50 343597 62 344573
rect 96 343597 108 344573
rect 50 343585 108 343597
rect -108 343355 -50 343367
rect -108 342379 -96 343355
rect -62 342379 -50 343355
rect -108 342367 -50 342379
rect 50 343355 108 343367
rect 50 342379 62 343355
rect 96 342379 108 343355
rect 50 342367 108 342379
rect -108 342137 -50 342149
rect -108 341161 -96 342137
rect -62 341161 -50 342137
rect -108 341149 -50 341161
rect 50 342137 108 342149
rect 50 341161 62 342137
rect 96 341161 108 342137
rect 50 341149 108 341161
rect -108 340919 -50 340931
rect -108 339943 -96 340919
rect -62 339943 -50 340919
rect -108 339931 -50 339943
rect 50 340919 108 340931
rect 50 339943 62 340919
rect 96 339943 108 340919
rect 50 339931 108 339943
rect -108 339701 -50 339713
rect -108 338725 -96 339701
rect -62 338725 -50 339701
rect -108 338713 -50 338725
rect 50 339701 108 339713
rect 50 338725 62 339701
rect 96 338725 108 339701
rect 50 338713 108 338725
rect -108 338483 -50 338495
rect -108 337507 -96 338483
rect -62 337507 -50 338483
rect -108 337495 -50 337507
rect 50 338483 108 338495
rect 50 337507 62 338483
rect 96 337507 108 338483
rect 50 337495 108 337507
rect -108 337265 -50 337277
rect -108 336289 -96 337265
rect -62 336289 -50 337265
rect -108 336277 -50 336289
rect 50 337265 108 337277
rect 50 336289 62 337265
rect 96 336289 108 337265
rect 50 336277 108 336289
rect -108 336047 -50 336059
rect -108 335071 -96 336047
rect -62 335071 -50 336047
rect -108 335059 -50 335071
rect 50 336047 108 336059
rect 50 335071 62 336047
rect 96 335071 108 336047
rect 50 335059 108 335071
rect -108 334829 -50 334841
rect -108 333853 -96 334829
rect -62 333853 -50 334829
rect -108 333841 -50 333853
rect 50 334829 108 334841
rect 50 333853 62 334829
rect 96 333853 108 334829
rect 50 333841 108 333853
rect -108 333611 -50 333623
rect -108 332635 -96 333611
rect -62 332635 -50 333611
rect -108 332623 -50 332635
rect 50 333611 108 333623
rect 50 332635 62 333611
rect 96 332635 108 333611
rect 50 332623 108 332635
rect -108 332393 -50 332405
rect -108 331417 -96 332393
rect -62 331417 -50 332393
rect -108 331405 -50 331417
rect 50 332393 108 332405
rect 50 331417 62 332393
rect 96 331417 108 332393
rect 50 331405 108 331417
rect -108 331175 -50 331187
rect -108 330199 -96 331175
rect -62 330199 -50 331175
rect -108 330187 -50 330199
rect 50 331175 108 331187
rect 50 330199 62 331175
rect 96 330199 108 331175
rect 50 330187 108 330199
rect -108 329957 -50 329969
rect -108 328981 -96 329957
rect -62 328981 -50 329957
rect -108 328969 -50 328981
rect 50 329957 108 329969
rect 50 328981 62 329957
rect 96 328981 108 329957
rect 50 328969 108 328981
rect -108 328739 -50 328751
rect -108 327763 -96 328739
rect -62 327763 -50 328739
rect -108 327751 -50 327763
rect 50 328739 108 328751
rect 50 327763 62 328739
rect 96 327763 108 328739
rect 50 327751 108 327763
rect -108 327521 -50 327533
rect -108 326545 -96 327521
rect -62 326545 -50 327521
rect -108 326533 -50 326545
rect 50 327521 108 327533
rect 50 326545 62 327521
rect 96 326545 108 327521
rect 50 326533 108 326545
rect -108 326303 -50 326315
rect -108 325327 -96 326303
rect -62 325327 -50 326303
rect -108 325315 -50 325327
rect 50 326303 108 326315
rect 50 325327 62 326303
rect 96 325327 108 326303
rect 50 325315 108 325327
rect -108 325085 -50 325097
rect -108 324109 -96 325085
rect -62 324109 -50 325085
rect -108 324097 -50 324109
rect 50 325085 108 325097
rect 50 324109 62 325085
rect 96 324109 108 325085
rect 50 324097 108 324109
rect -108 323867 -50 323879
rect -108 322891 -96 323867
rect -62 322891 -50 323867
rect -108 322879 -50 322891
rect 50 323867 108 323879
rect 50 322891 62 323867
rect 96 322891 108 323867
rect 50 322879 108 322891
rect -108 322649 -50 322661
rect -108 321673 -96 322649
rect -62 321673 -50 322649
rect -108 321661 -50 321673
rect 50 322649 108 322661
rect 50 321673 62 322649
rect 96 321673 108 322649
rect 50 321661 108 321673
rect -108 321431 -50 321443
rect -108 320455 -96 321431
rect -62 320455 -50 321431
rect -108 320443 -50 320455
rect 50 321431 108 321443
rect 50 320455 62 321431
rect 96 320455 108 321431
rect 50 320443 108 320455
rect -108 320213 -50 320225
rect -108 319237 -96 320213
rect -62 319237 -50 320213
rect -108 319225 -50 319237
rect 50 320213 108 320225
rect 50 319237 62 320213
rect 96 319237 108 320213
rect 50 319225 108 319237
rect -108 318995 -50 319007
rect -108 318019 -96 318995
rect -62 318019 -50 318995
rect -108 318007 -50 318019
rect 50 318995 108 319007
rect 50 318019 62 318995
rect 96 318019 108 318995
rect 50 318007 108 318019
rect -108 317777 -50 317789
rect -108 316801 -96 317777
rect -62 316801 -50 317777
rect -108 316789 -50 316801
rect 50 317777 108 317789
rect 50 316801 62 317777
rect 96 316801 108 317777
rect 50 316789 108 316801
rect -108 316559 -50 316571
rect -108 315583 -96 316559
rect -62 315583 -50 316559
rect -108 315571 -50 315583
rect 50 316559 108 316571
rect 50 315583 62 316559
rect 96 315583 108 316559
rect 50 315571 108 315583
rect -108 315341 -50 315353
rect -108 314365 -96 315341
rect -62 314365 -50 315341
rect -108 314353 -50 314365
rect 50 315341 108 315353
rect 50 314365 62 315341
rect 96 314365 108 315341
rect 50 314353 108 314365
rect -108 314123 -50 314135
rect -108 313147 -96 314123
rect -62 313147 -50 314123
rect -108 313135 -50 313147
rect 50 314123 108 314135
rect 50 313147 62 314123
rect 96 313147 108 314123
rect 50 313135 108 313147
rect -108 312905 -50 312917
rect -108 311929 -96 312905
rect -62 311929 -50 312905
rect -108 311917 -50 311929
rect 50 312905 108 312917
rect 50 311929 62 312905
rect 96 311929 108 312905
rect 50 311917 108 311929
rect -108 311687 -50 311699
rect -108 310711 -96 311687
rect -62 310711 -50 311687
rect -108 310699 -50 310711
rect 50 311687 108 311699
rect 50 310711 62 311687
rect 96 310711 108 311687
rect 50 310699 108 310711
rect -108 310469 -50 310481
rect -108 309493 -96 310469
rect -62 309493 -50 310469
rect -108 309481 -50 309493
rect 50 310469 108 310481
rect 50 309493 62 310469
rect 96 309493 108 310469
rect 50 309481 108 309493
rect -108 309251 -50 309263
rect -108 308275 -96 309251
rect -62 308275 -50 309251
rect -108 308263 -50 308275
rect 50 309251 108 309263
rect 50 308275 62 309251
rect 96 308275 108 309251
rect 50 308263 108 308275
rect -108 308033 -50 308045
rect -108 307057 -96 308033
rect -62 307057 -50 308033
rect -108 307045 -50 307057
rect 50 308033 108 308045
rect 50 307057 62 308033
rect 96 307057 108 308033
rect 50 307045 108 307057
rect -108 306815 -50 306827
rect -108 305839 -96 306815
rect -62 305839 -50 306815
rect -108 305827 -50 305839
rect 50 306815 108 306827
rect 50 305839 62 306815
rect 96 305839 108 306815
rect 50 305827 108 305839
rect -108 305597 -50 305609
rect -108 304621 -96 305597
rect -62 304621 -50 305597
rect -108 304609 -50 304621
rect 50 305597 108 305609
rect 50 304621 62 305597
rect 96 304621 108 305597
rect 50 304609 108 304621
rect -108 304379 -50 304391
rect -108 303403 -96 304379
rect -62 303403 -50 304379
rect -108 303391 -50 303403
rect 50 304379 108 304391
rect 50 303403 62 304379
rect 96 303403 108 304379
rect 50 303391 108 303403
rect -108 303161 -50 303173
rect -108 302185 -96 303161
rect -62 302185 -50 303161
rect -108 302173 -50 302185
rect 50 303161 108 303173
rect 50 302185 62 303161
rect 96 302185 108 303161
rect 50 302173 108 302185
rect -108 301943 -50 301955
rect -108 300967 -96 301943
rect -62 300967 -50 301943
rect -108 300955 -50 300967
rect 50 301943 108 301955
rect 50 300967 62 301943
rect 96 300967 108 301943
rect 50 300955 108 300967
rect -108 300725 -50 300737
rect -108 299749 -96 300725
rect -62 299749 -50 300725
rect -108 299737 -50 299749
rect 50 300725 108 300737
rect 50 299749 62 300725
rect 96 299749 108 300725
rect 50 299737 108 299749
rect -108 299507 -50 299519
rect -108 298531 -96 299507
rect -62 298531 -50 299507
rect -108 298519 -50 298531
rect 50 299507 108 299519
rect 50 298531 62 299507
rect 96 298531 108 299507
rect 50 298519 108 298531
rect -108 298289 -50 298301
rect -108 297313 -96 298289
rect -62 297313 -50 298289
rect -108 297301 -50 297313
rect 50 298289 108 298301
rect 50 297313 62 298289
rect 96 297313 108 298289
rect 50 297301 108 297313
rect -108 297071 -50 297083
rect -108 296095 -96 297071
rect -62 296095 -50 297071
rect -108 296083 -50 296095
rect 50 297071 108 297083
rect 50 296095 62 297071
rect 96 296095 108 297071
rect 50 296083 108 296095
rect -108 295853 -50 295865
rect -108 294877 -96 295853
rect -62 294877 -50 295853
rect -108 294865 -50 294877
rect 50 295853 108 295865
rect 50 294877 62 295853
rect 96 294877 108 295853
rect 50 294865 108 294877
rect -108 294635 -50 294647
rect -108 293659 -96 294635
rect -62 293659 -50 294635
rect -108 293647 -50 293659
rect 50 294635 108 294647
rect 50 293659 62 294635
rect 96 293659 108 294635
rect 50 293647 108 293659
rect -108 293417 -50 293429
rect -108 292441 -96 293417
rect -62 292441 -50 293417
rect -108 292429 -50 292441
rect 50 293417 108 293429
rect 50 292441 62 293417
rect 96 292441 108 293417
rect 50 292429 108 292441
rect -108 292199 -50 292211
rect -108 291223 -96 292199
rect -62 291223 -50 292199
rect -108 291211 -50 291223
rect 50 292199 108 292211
rect 50 291223 62 292199
rect 96 291223 108 292199
rect 50 291211 108 291223
rect -108 290981 -50 290993
rect -108 290005 -96 290981
rect -62 290005 -50 290981
rect -108 289993 -50 290005
rect 50 290981 108 290993
rect 50 290005 62 290981
rect 96 290005 108 290981
rect 50 289993 108 290005
rect -108 289763 -50 289775
rect -108 288787 -96 289763
rect -62 288787 -50 289763
rect -108 288775 -50 288787
rect 50 289763 108 289775
rect 50 288787 62 289763
rect 96 288787 108 289763
rect 50 288775 108 288787
rect -108 288545 -50 288557
rect -108 287569 -96 288545
rect -62 287569 -50 288545
rect -108 287557 -50 287569
rect 50 288545 108 288557
rect 50 287569 62 288545
rect 96 287569 108 288545
rect 50 287557 108 287569
rect -108 287327 -50 287339
rect -108 286351 -96 287327
rect -62 286351 -50 287327
rect -108 286339 -50 286351
rect 50 287327 108 287339
rect 50 286351 62 287327
rect 96 286351 108 287327
rect 50 286339 108 286351
rect -108 286109 -50 286121
rect -108 285133 -96 286109
rect -62 285133 -50 286109
rect -108 285121 -50 285133
rect 50 286109 108 286121
rect 50 285133 62 286109
rect 96 285133 108 286109
rect 50 285121 108 285133
rect -108 284891 -50 284903
rect -108 283915 -96 284891
rect -62 283915 -50 284891
rect -108 283903 -50 283915
rect 50 284891 108 284903
rect 50 283915 62 284891
rect 96 283915 108 284891
rect 50 283903 108 283915
rect -108 283673 -50 283685
rect -108 282697 -96 283673
rect -62 282697 -50 283673
rect -108 282685 -50 282697
rect 50 283673 108 283685
rect 50 282697 62 283673
rect 96 282697 108 283673
rect 50 282685 108 282697
rect -108 282455 -50 282467
rect -108 281479 -96 282455
rect -62 281479 -50 282455
rect -108 281467 -50 281479
rect 50 282455 108 282467
rect 50 281479 62 282455
rect 96 281479 108 282455
rect 50 281467 108 281479
rect -108 281237 -50 281249
rect -108 280261 -96 281237
rect -62 280261 -50 281237
rect -108 280249 -50 280261
rect 50 281237 108 281249
rect 50 280261 62 281237
rect 96 280261 108 281237
rect 50 280249 108 280261
rect -108 280019 -50 280031
rect -108 279043 -96 280019
rect -62 279043 -50 280019
rect -108 279031 -50 279043
rect 50 280019 108 280031
rect 50 279043 62 280019
rect 96 279043 108 280019
rect 50 279031 108 279043
rect -108 278801 -50 278813
rect -108 277825 -96 278801
rect -62 277825 -50 278801
rect -108 277813 -50 277825
rect 50 278801 108 278813
rect 50 277825 62 278801
rect 96 277825 108 278801
rect 50 277813 108 277825
rect -108 277583 -50 277595
rect -108 276607 -96 277583
rect -62 276607 -50 277583
rect -108 276595 -50 276607
rect 50 277583 108 277595
rect 50 276607 62 277583
rect 96 276607 108 277583
rect 50 276595 108 276607
rect -108 276365 -50 276377
rect -108 275389 -96 276365
rect -62 275389 -50 276365
rect -108 275377 -50 275389
rect 50 276365 108 276377
rect 50 275389 62 276365
rect 96 275389 108 276365
rect 50 275377 108 275389
rect -108 275147 -50 275159
rect -108 274171 -96 275147
rect -62 274171 -50 275147
rect -108 274159 -50 274171
rect 50 275147 108 275159
rect 50 274171 62 275147
rect 96 274171 108 275147
rect 50 274159 108 274171
rect -108 273929 -50 273941
rect -108 272953 -96 273929
rect -62 272953 -50 273929
rect -108 272941 -50 272953
rect 50 273929 108 273941
rect 50 272953 62 273929
rect 96 272953 108 273929
rect 50 272941 108 272953
rect -108 272711 -50 272723
rect -108 271735 -96 272711
rect -62 271735 -50 272711
rect -108 271723 -50 271735
rect 50 272711 108 272723
rect 50 271735 62 272711
rect 96 271735 108 272711
rect 50 271723 108 271735
rect -108 271493 -50 271505
rect -108 270517 -96 271493
rect -62 270517 -50 271493
rect -108 270505 -50 270517
rect 50 271493 108 271505
rect 50 270517 62 271493
rect 96 270517 108 271493
rect 50 270505 108 270517
rect -108 270275 -50 270287
rect -108 269299 -96 270275
rect -62 269299 -50 270275
rect -108 269287 -50 269299
rect 50 270275 108 270287
rect 50 269299 62 270275
rect 96 269299 108 270275
rect 50 269287 108 269299
rect -108 269057 -50 269069
rect -108 268081 -96 269057
rect -62 268081 -50 269057
rect -108 268069 -50 268081
rect 50 269057 108 269069
rect 50 268081 62 269057
rect 96 268081 108 269057
rect 50 268069 108 268081
rect -108 267839 -50 267851
rect -108 266863 -96 267839
rect -62 266863 -50 267839
rect -108 266851 -50 266863
rect 50 267839 108 267851
rect 50 266863 62 267839
rect 96 266863 108 267839
rect 50 266851 108 266863
rect -108 266621 -50 266633
rect -108 265645 -96 266621
rect -62 265645 -50 266621
rect -108 265633 -50 265645
rect 50 266621 108 266633
rect 50 265645 62 266621
rect 96 265645 108 266621
rect 50 265633 108 265645
rect -108 265403 -50 265415
rect -108 264427 -96 265403
rect -62 264427 -50 265403
rect -108 264415 -50 264427
rect 50 265403 108 265415
rect 50 264427 62 265403
rect 96 264427 108 265403
rect 50 264415 108 264427
rect -108 264185 -50 264197
rect -108 263209 -96 264185
rect -62 263209 -50 264185
rect -108 263197 -50 263209
rect 50 264185 108 264197
rect 50 263209 62 264185
rect 96 263209 108 264185
rect 50 263197 108 263209
rect -108 262967 -50 262979
rect -108 261991 -96 262967
rect -62 261991 -50 262967
rect -108 261979 -50 261991
rect 50 262967 108 262979
rect 50 261991 62 262967
rect 96 261991 108 262967
rect 50 261979 108 261991
rect -108 261749 -50 261761
rect -108 260773 -96 261749
rect -62 260773 -50 261749
rect -108 260761 -50 260773
rect 50 261749 108 261761
rect 50 260773 62 261749
rect 96 260773 108 261749
rect 50 260761 108 260773
rect -108 260531 -50 260543
rect -108 259555 -96 260531
rect -62 259555 -50 260531
rect -108 259543 -50 259555
rect 50 260531 108 260543
rect 50 259555 62 260531
rect 96 259555 108 260531
rect 50 259543 108 259555
rect -108 259313 -50 259325
rect -108 258337 -96 259313
rect -62 258337 -50 259313
rect -108 258325 -50 258337
rect 50 259313 108 259325
rect 50 258337 62 259313
rect 96 258337 108 259313
rect 50 258325 108 258337
rect -108 258095 -50 258107
rect -108 257119 -96 258095
rect -62 257119 -50 258095
rect -108 257107 -50 257119
rect 50 258095 108 258107
rect 50 257119 62 258095
rect 96 257119 108 258095
rect 50 257107 108 257119
rect -108 256877 -50 256889
rect -108 255901 -96 256877
rect -62 255901 -50 256877
rect -108 255889 -50 255901
rect 50 256877 108 256889
rect 50 255901 62 256877
rect 96 255901 108 256877
rect 50 255889 108 255901
rect -108 255659 -50 255671
rect -108 254683 -96 255659
rect -62 254683 -50 255659
rect -108 254671 -50 254683
rect 50 255659 108 255671
rect 50 254683 62 255659
rect 96 254683 108 255659
rect 50 254671 108 254683
rect -108 254441 -50 254453
rect -108 253465 -96 254441
rect -62 253465 -50 254441
rect -108 253453 -50 253465
rect 50 254441 108 254453
rect 50 253465 62 254441
rect 96 253465 108 254441
rect 50 253453 108 253465
rect -108 253223 -50 253235
rect -108 252247 -96 253223
rect -62 252247 -50 253223
rect -108 252235 -50 252247
rect 50 253223 108 253235
rect 50 252247 62 253223
rect 96 252247 108 253223
rect 50 252235 108 252247
rect -108 252005 -50 252017
rect -108 251029 -96 252005
rect -62 251029 -50 252005
rect -108 251017 -50 251029
rect 50 252005 108 252017
rect 50 251029 62 252005
rect 96 251029 108 252005
rect 50 251017 108 251029
rect -108 250787 -50 250799
rect -108 249811 -96 250787
rect -62 249811 -50 250787
rect -108 249799 -50 249811
rect 50 250787 108 250799
rect 50 249811 62 250787
rect 96 249811 108 250787
rect 50 249799 108 249811
rect -108 249569 -50 249581
rect -108 248593 -96 249569
rect -62 248593 -50 249569
rect -108 248581 -50 248593
rect 50 249569 108 249581
rect 50 248593 62 249569
rect 96 248593 108 249569
rect 50 248581 108 248593
rect -108 248351 -50 248363
rect -108 247375 -96 248351
rect -62 247375 -50 248351
rect -108 247363 -50 247375
rect 50 248351 108 248363
rect 50 247375 62 248351
rect 96 247375 108 248351
rect 50 247363 108 247375
rect -108 247133 -50 247145
rect -108 246157 -96 247133
rect -62 246157 -50 247133
rect -108 246145 -50 246157
rect 50 247133 108 247145
rect 50 246157 62 247133
rect 96 246157 108 247133
rect 50 246145 108 246157
rect -108 245915 -50 245927
rect -108 244939 -96 245915
rect -62 244939 -50 245915
rect -108 244927 -50 244939
rect 50 245915 108 245927
rect 50 244939 62 245915
rect 96 244939 108 245915
rect 50 244927 108 244939
rect -108 244697 -50 244709
rect -108 243721 -96 244697
rect -62 243721 -50 244697
rect -108 243709 -50 243721
rect 50 244697 108 244709
rect 50 243721 62 244697
rect 96 243721 108 244697
rect 50 243709 108 243721
rect -108 243479 -50 243491
rect -108 242503 -96 243479
rect -62 242503 -50 243479
rect -108 242491 -50 242503
rect 50 243479 108 243491
rect 50 242503 62 243479
rect 96 242503 108 243479
rect 50 242491 108 242503
rect -108 242261 -50 242273
rect -108 241285 -96 242261
rect -62 241285 -50 242261
rect -108 241273 -50 241285
rect 50 242261 108 242273
rect 50 241285 62 242261
rect 96 241285 108 242261
rect 50 241273 108 241285
rect -108 241043 -50 241055
rect -108 240067 -96 241043
rect -62 240067 -50 241043
rect -108 240055 -50 240067
rect 50 241043 108 241055
rect 50 240067 62 241043
rect 96 240067 108 241043
rect 50 240055 108 240067
rect -108 239825 -50 239837
rect -108 238849 -96 239825
rect -62 238849 -50 239825
rect -108 238837 -50 238849
rect 50 239825 108 239837
rect 50 238849 62 239825
rect 96 238849 108 239825
rect 50 238837 108 238849
rect -108 238607 -50 238619
rect -108 237631 -96 238607
rect -62 237631 -50 238607
rect -108 237619 -50 237631
rect 50 238607 108 238619
rect 50 237631 62 238607
rect 96 237631 108 238607
rect 50 237619 108 237631
rect -108 237389 -50 237401
rect -108 236413 -96 237389
rect -62 236413 -50 237389
rect -108 236401 -50 236413
rect 50 237389 108 237401
rect 50 236413 62 237389
rect 96 236413 108 237389
rect 50 236401 108 236413
rect -108 236171 -50 236183
rect -108 235195 -96 236171
rect -62 235195 -50 236171
rect -108 235183 -50 235195
rect 50 236171 108 236183
rect 50 235195 62 236171
rect 96 235195 108 236171
rect 50 235183 108 235195
rect -108 234953 -50 234965
rect -108 233977 -96 234953
rect -62 233977 -50 234953
rect -108 233965 -50 233977
rect 50 234953 108 234965
rect 50 233977 62 234953
rect 96 233977 108 234953
rect 50 233965 108 233977
rect -108 233735 -50 233747
rect -108 232759 -96 233735
rect -62 232759 -50 233735
rect -108 232747 -50 232759
rect 50 233735 108 233747
rect 50 232759 62 233735
rect 96 232759 108 233735
rect 50 232747 108 232759
rect -108 232517 -50 232529
rect -108 231541 -96 232517
rect -62 231541 -50 232517
rect -108 231529 -50 231541
rect 50 232517 108 232529
rect 50 231541 62 232517
rect 96 231541 108 232517
rect 50 231529 108 231541
rect -108 231299 -50 231311
rect -108 230323 -96 231299
rect -62 230323 -50 231299
rect -108 230311 -50 230323
rect 50 231299 108 231311
rect 50 230323 62 231299
rect 96 230323 108 231299
rect 50 230311 108 230323
rect -108 230081 -50 230093
rect -108 229105 -96 230081
rect -62 229105 -50 230081
rect -108 229093 -50 229105
rect 50 230081 108 230093
rect 50 229105 62 230081
rect 96 229105 108 230081
rect 50 229093 108 229105
rect -108 228863 -50 228875
rect -108 227887 -96 228863
rect -62 227887 -50 228863
rect -108 227875 -50 227887
rect 50 228863 108 228875
rect 50 227887 62 228863
rect 96 227887 108 228863
rect 50 227875 108 227887
rect -108 227645 -50 227657
rect -108 226669 -96 227645
rect -62 226669 -50 227645
rect -108 226657 -50 226669
rect 50 227645 108 227657
rect 50 226669 62 227645
rect 96 226669 108 227645
rect 50 226657 108 226669
rect -108 226427 -50 226439
rect -108 225451 -96 226427
rect -62 225451 -50 226427
rect -108 225439 -50 225451
rect 50 226427 108 226439
rect 50 225451 62 226427
rect 96 225451 108 226427
rect 50 225439 108 225451
rect -108 225209 -50 225221
rect -108 224233 -96 225209
rect -62 224233 -50 225209
rect -108 224221 -50 224233
rect 50 225209 108 225221
rect 50 224233 62 225209
rect 96 224233 108 225209
rect 50 224221 108 224233
rect -108 223991 -50 224003
rect -108 223015 -96 223991
rect -62 223015 -50 223991
rect -108 223003 -50 223015
rect 50 223991 108 224003
rect 50 223015 62 223991
rect 96 223015 108 223991
rect 50 223003 108 223015
rect -108 222773 -50 222785
rect -108 221797 -96 222773
rect -62 221797 -50 222773
rect -108 221785 -50 221797
rect 50 222773 108 222785
rect 50 221797 62 222773
rect 96 221797 108 222773
rect 50 221785 108 221797
rect -108 221555 -50 221567
rect -108 220579 -96 221555
rect -62 220579 -50 221555
rect -108 220567 -50 220579
rect 50 221555 108 221567
rect 50 220579 62 221555
rect 96 220579 108 221555
rect 50 220567 108 220579
rect -108 220337 -50 220349
rect -108 219361 -96 220337
rect -62 219361 -50 220337
rect -108 219349 -50 219361
rect 50 220337 108 220349
rect 50 219361 62 220337
rect 96 219361 108 220337
rect 50 219349 108 219361
rect -108 219119 -50 219131
rect -108 218143 -96 219119
rect -62 218143 -50 219119
rect -108 218131 -50 218143
rect 50 219119 108 219131
rect 50 218143 62 219119
rect 96 218143 108 219119
rect 50 218131 108 218143
rect -108 217901 -50 217913
rect -108 216925 -96 217901
rect -62 216925 -50 217901
rect -108 216913 -50 216925
rect 50 217901 108 217913
rect 50 216925 62 217901
rect 96 216925 108 217901
rect 50 216913 108 216925
rect -108 216683 -50 216695
rect -108 215707 -96 216683
rect -62 215707 -50 216683
rect -108 215695 -50 215707
rect 50 216683 108 216695
rect 50 215707 62 216683
rect 96 215707 108 216683
rect 50 215695 108 215707
rect -108 215465 -50 215477
rect -108 214489 -96 215465
rect -62 214489 -50 215465
rect -108 214477 -50 214489
rect 50 215465 108 215477
rect 50 214489 62 215465
rect 96 214489 108 215465
rect 50 214477 108 214489
rect -108 214247 -50 214259
rect -108 213271 -96 214247
rect -62 213271 -50 214247
rect -108 213259 -50 213271
rect 50 214247 108 214259
rect 50 213271 62 214247
rect 96 213271 108 214247
rect 50 213259 108 213271
rect -108 213029 -50 213041
rect -108 212053 -96 213029
rect -62 212053 -50 213029
rect -108 212041 -50 212053
rect 50 213029 108 213041
rect 50 212053 62 213029
rect 96 212053 108 213029
rect 50 212041 108 212053
rect -108 211811 -50 211823
rect -108 210835 -96 211811
rect -62 210835 -50 211811
rect -108 210823 -50 210835
rect 50 211811 108 211823
rect 50 210835 62 211811
rect 96 210835 108 211811
rect 50 210823 108 210835
rect -108 210593 -50 210605
rect -108 209617 -96 210593
rect -62 209617 -50 210593
rect -108 209605 -50 209617
rect 50 210593 108 210605
rect 50 209617 62 210593
rect 96 209617 108 210593
rect 50 209605 108 209617
rect -108 209375 -50 209387
rect -108 208399 -96 209375
rect -62 208399 -50 209375
rect -108 208387 -50 208399
rect 50 209375 108 209387
rect 50 208399 62 209375
rect 96 208399 108 209375
rect 50 208387 108 208399
rect -108 208157 -50 208169
rect -108 207181 -96 208157
rect -62 207181 -50 208157
rect -108 207169 -50 207181
rect 50 208157 108 208169
rect 50 207181 62 208157
rect 96 207181 108 208157
rect 50 207169 108 207181
rect -108 206939 -50 206951
rect -108 205963 -96 206939
rect -62 205963 -50 206939
rect -108 205951 -50 205963
rect 50 206939 108 206951
rect 50 205963 62 206939
rect 96 205963 108 206939
rect 50 205951 108 205963
rect -108 205721 -50 205733
rect -108 204745 -96 205721
rect -62 204745 -50 205721
rect -108 204733 -50 204745
rect 50 205721 108 205733
rect 50 204745 62 205721
rect 96 204745 108 205721
rect 50 204733 108 204745
rect -108 204503 -50 204515
rect -108 203527 -96 204503
rect -62 203527 -50 204503
rect -108 203515 -50 203527
rect 50 204503 108 204515
rect 50 203527 62 204503
rect 96 203527 108 204503
rect 50 203515 108 203527
rect -108 203285 -50 203297
rect -108 202309 -96 203285
rect -62 202309 -50 203285
rect -108 202297 -50 202309
rect 50 203285 108 203297
rect 50 202309 62 203285
rect 96 202309 108 203285
rect 50 202297 108 202309
rect -108 202067 -50 202079
rect -108 201091 -96 202067
rect -62 201091 -50 202067
rect -108 201079 -50 201091
rect 50 202067 108 202079
rect 50 201091 62 202067
rect 96 201091 108 202067
rect 50 201079 108 201091
rect -108 200849 -50 200861
rect -108 199873 -96 200849
rect -62 199873 -50 200849
rect -108 199861 -50 199873
rect 50 200849 108 200861
rect 50 199873 62 200849
rect 96 199873 108 200849
rect 50 199861 108 199873
rect -108 199631 -50 199643
rect -108 198655 -96 199631
rect -62 198655 -50 199631
rect -108 198643 -50 198655
rect 50 199631 108 199643
rect 50 198655 62 199631
rect 96 198655 108 199631
rect 50 198643 108 198655
rect -108 198413 -50 198425
rect -108 197437 -96 198413
rect -62 197437 -50 198413
rect -108 197425 -50 197437
rect 50 198413 108 198425
rect 50 197437 62 198413
rect 96 197437 108 198413
rect 50 197425 108 197437
rect -108 197195 -50 197207
rect -108 196219 -96 197195
rect -62 196219 -50 197195
rect -108 196207 -50 196219
rect 50 197195 108 197207
rect 50 196219 62 197195
rect 96 196219 108 197195
rect 50 196207 108 196219
rect -108 195977 -50 195989
rect -108 195001 -96 195977
rect -62 195001 -50 195977
rect -108 194989 -50 195001
rect 50 195977 108 195989
rect 50 195001 62 195977
rect 96 195001 108 195977
rect 50 194989 108 195001
rect -108 194759 -50 194771
rect -108 193783 -96 194759
rect -62 193783 -50 194759
rect -108 193771 -50 193783
rect 50 194759 108 194771
rect 50 193783 62 194759
rect 96 193783 108 194759
rect 50 193771 108 193783
rect -108 193541 -50 193553
rect -108 192565 -96 193541
rect -62 192565 -50 193541
rect -108 192553 -50 192565
rect 50 193541 108 193553
rect 50 192565 62 193541
rect 96 192565 108 193541
rect 50 192553 108 192565
rect -108 192323 -50 192335
rect -108 191347 -96 192323
rect -62 191347 -50 192323
rect -108 191335 -50 191347
rect 50 192323 108 192335
rect 50 191347 62 192323
rect 96 191347 108 192323
rect 50 191335 108 191347
rect -108 191105 -50 191117
rect -108 190129 -96 191105
rect -62 190129 -50 191105
rect -108 190117 -50 190129
rect 50 191105 108 191117
rect 50 190129 62 191105
rect 96 190129 108 191105
rect 50 190117 108 190129
rect -108 189887 -50 189899
rect -108 188911 -96 189887
rect -62 188911 -50 189887
rect -108 188899 -50 188911
rect 50 189887 108 189899
rect 50 188911 62 189887
rect 96 188911 108 189887
rect 50 188899 108 188911
rect -108 188669 -50 188681
rect -108 187693 -96 188669
rect -62 187693 -50 188669
rect -108 187681 -50 187693
rect 50 188669 108 188681
rect 50 187693 62 188669
rect 96 187693 108 188669
rect 50 187681 108 187693
rect -108 187451 -50 187463
rect -108 186475 -96 187451
rect -62 186475 -50 187451
rect -108 186463 -50 186475
rect 50 187451 108 187463
rect 50 186475 62 187451
rect 96 186475 108 187451
rect 50 186463 108 186475
rect -108 186233 -50 186245
rect -108 185257 -96 186233
rect -62 185257 -50 186233
rect -108 185245 -50 185257
rect 50 186233 108 186245
rect 50 185257 62 186233
rect 96 185257 108 186233
rect 50 185245 108 185257
rect -108 185015 -50 185027
rect -108 184039 -96 185015
rect -62 184039 -50 185015
rect -108 184027 -50 184039
rect 50 185015 108 185027
rect 50 184039 62 185015
rect 96 184039 108 185015
rect 50 184027 108 184039
rect -108 183797 -50 183809
rect -108 182821 -96 183797
rect -62 182821 -50 183797
rect -108 182809 -50 182821
rect 50 183797 108 183809
rect 50 182821 62 183797
rect 96 182821 108 183797
rect 50 182809 108 182821
rect -108 182579 -50 182591
rect -108 181603 -96 182579
rect -62 181603 -50 182579
rect -108 181591 -50 181603
rect 50 182579 108 182591
rect 50 181603 62 182579
rect 96 181603 108 182579
rect 50 181591 108 181603
rect -108 181361 -50 181373
rect -108 180385 -96 181361
rect -62 180385 -50 181361
rect -108 180373 -50 180385
rect 50 181361 108 181373
rect 50 180385 62 181361
rect 96 180385 108 181361
rect 50 180373 108 180385
rect -108 180143 -50 180155
rect -108 179167 -96 180143
rect -62 179167 -50 180143
rect -108 179155 -50 179167
rect 50 180143 108 180155
rect 50 179167 62 180143
rect 96 179167 108 180143
rect 50 179155 108 179167
rect -108 178925 -50 178937
rect -108 177949 -96 178925
rect -62 177949 -50 178925
rect -108 177937 -50 177949
rect 50 178925 108 178937
rect 50 177949 62 178925
rect 96 177949 108 178925
rect 50 177937 108 177949
rect -108 177707 -50 177719
rect -108 176731 -96 177707
rect -62 176731 -50 177707
rect -108 176719 -50 176731
rect 50 177707 108 177719
rect 50 176731 62 177707
rect 96 176731 108 177707
rect 50 176719 108 176731
rect -108 176489 -50 176501
rect -108 175513 -96 176489
rect -62 175513 -50 176489
rect -108 175501 -50 175513
rect 50 176489 108 176501
rect 50 175513 62 176489
rect 96 175513 108 176489
rect 50 175501 108 175513
rect -108 175271 -50 175283
rect -108 174295 -96 175271
rect -62 174295 -50 175271
rect -108 174283 -50 174295
rect 50 175271 108 175283
rect 50 174295 62 175271
rect 96 174295 108 175271
rect 50 174283 108 174295
rect -108 174053 -50 174065
rect -108 173077 -96 174053
rect -62 173077 -50 174053
rect -108 173065 -50 173077
rect 50 174053 108 174065
rect 50 173077 62 174053
rect 96 173077 108 174053
rect 50 173065 108 173077
rect -108 172835 -50 172847
rect -108 171859 -96 172835
rect -62 171859 -50 172835
rect -108 171847 -50 171859
rect 50 172835 108 172847
rect 50 171859 62 172835
rect 96 171859 108 172835
rect 50 171847 108 171859
rect -108 171617 -50 171629
rect -108 170641 -96 171617
rect -62 170641 -50 171617
rect -108 170629 -50 170641
rect 50 171617 108 171629
rect 50 170641 62 171617
rect 96 170641 108 171617
rect 50 170629 108 170641
rect -108 170399 -50 170411
rect -108 169423 -96 170399
rect -62 169423 -50 170399
rect -108 169411 -50 169423
rect 50 170399 108 170411
rect 50 169423 62 170399
rect 96 169423 108 170399
rect 50 169411 108 169423
rect -108 169181 -50 169193
rect -108 168205 -96 169181
rect -62 168205 -50 169181
rect -108 168193 -50 168205
rect 50 169181 108 169193
rect 50 168205 62 169181
rect 96 168205 108 169181
rect 50 168193 108 168205
rect -108 167963 -50 167975
rect -108 166987 -96 167963
rect -62 166987 -50 167963
rect -108 166975 -50 166987
rect 50 167963 108 167975
rect 50 166987 62 167963
rect 96 166987 108 167963
rect 50 166975 108 166987
rect -108 166745 -50 166757
rect -108 165769 -96 166745
rect -62 165769 -50 166745
rect -108 165757 -50 165769
rect 50 166745 108 166757
rect 50 165769 62 166745
rect 96 165769 108 166745
rect 50 165757 108 165769
rect -108 165527 -50 165539
rect -108 164551 -96 165527
rect -62 164551 -50 165527
rect -108 164539 -50 164551
rect 50 165527 108 165539
rect 50 164551 62 165527
rect 96 164551 108 165527
rect 50 164539 108 164551
rect -108 164309 -50 164321
rect -108 163333 -96 164309
rect -62 163333 -50 164309
rect -108 163321 -50 163333
rect 50 164309 108 164321
rect 50 163333 62 164309
rect 96 163333 108 164309
rect 50 163321 108 163333
rect -108 163091 -50 163103
rect -108 162115 -96 163091
rect -62 162115 -50 163091
rect -108 162103 -50 162115
rect 50 163091 108 163103
rect 50 162115 62 163091
rect 96 162115 108 163091
rect 50 162103 108 162115
rect -108 161873 -50 161885
rect -108 160897 -96 161873
rect -62 160897 -50 161873
rect -108 160885 -50 160897
rect 50 161873 108 161885
rect 50 160897 62 161873
rect 96 160897 108 161873
rect 50 160885 108 160897
rect -108 160655 -50 160667
rect -108 159679 -96 160655
rect -62 159679 -50 160655
rect -108 159667 -50 159679
rect 50 160655 108 160667
rect 50 159679 62 160655
rect 96 159679 108 160655
rect 50 159667 108 159679
rect -108 159437 -50 159449
rect -108 158461 -96 159437
rect -62 158461 -50 159437
rect -108 158449 -50 158461
rect 50 159437 108 159449
rect 50 158461 62 159437
rect 96 158461 108 159437
rect 50 158449 108 158461
rect -108 158219 -50 158231
rect -108 157243 -96 158219
rect -62 157243 -50 158219
rect -108 157231 -50 157243
rect 50 158219 108 158231
rect 50 157243 62 158219
rect 96 157243 108 158219
rect 50 157231 108 157243
rect -108 157001 -50 157013
rect -108 156025 -96 157001
rect -62 156025 -50 157001
rect -108 156013 -50 156025
rect 50 157001 108 157013
rect 50 156025 62 157001
rect 96 156025 108 157001
rect 50 156013 108 156025
rect -108 155783 -50 155795
rect -108 154807 -96 155783
rect -62 154807 -50 155783
rect -108 154795 -50 154807
rect 50 155783 108 155795
rect 50 154807 62 155783
rect 96 154807 108 155783
rect 50 154795 108 154807
rect -108 154565 -50 154577
rect -108 153589 -96 154565
rect -62 153589 -50 154565
rect -108 153577 -50 153589
rect 50 154565 108 154577
rect 50 153589 62 154565
rect 96 153589 108 154565
rect 50 153577 108 153589
rect -108 153347 -50 153359
rect -108 152371 -96 153347
rect -62 152371 -50 153347
rect -108 152359 -50 152371
rect 50 153347 108 153359
rect 50 152371 62 153347
rect 96 152371 108 153347
rect 50 152359 108 152371
rect -108 152129 -50 152141
rect -108 151153 -96 152129
rect -62 151153 -50 152129
rect -108 151141 -50 151153
rect 50 152129 108 152141
rect 50 151153 62 152129
rect 96 151153 108 152129
rect 50 151141 108 151153
rect -108 150911 -50 150923
rect -108 149935 -96 150911
rect -62 149935 -50 150911
rect -108 149923 -50 149935
rect 50 150911 108 150923
rect 50 149935 62 150911
rect 96 149935 108 150911
rect 50 149923 108 149935
rect -108 149693 -50 149705
rect -108 148717 -96 149693
rect -62 148717 -50 149693
rect -108 148705 -50 148717
rect 50 149693 108 149705
rect 50 148717 62 149693
rect 96 148717 108 149693
rect 50 148705 108 148717
rect -108 148475 -50 148487
rect -108 147499 -96 148475
rect -62 147499 -50 148475
rect -108 147487 -50 147499
rect 50 148475 108 148487
rect 50 147499 62 148475
rect 96 147499 108 148475
rect 50 147487 108 147499
rect -108 147257 -50 147269
rect -108 146281 -96 147257
rect -62 146281 -50 147257
rect -108 146269 -50 146281
rect 50 147257 108 147269
rect 50 146281 62 147257
rect 96 146281 108 147257
rect 50 146269 108 146281
rect -108 146039 -50 146051
rect -108 145063 -96 146039
rect -62 145063 -50 146039
rect -108 145051 -50 145063
rect 50 146039 108 146051
rect 50 145063 62 146039
rect 96 145063 108 146039
rect 50 145051 108 145063
rect -108 144821 -50 144833
rect -108 143845 -96 144821
rect -62 143845 -50 144821
rect -108 143833 -50 143845
rect 50 144821 108 144833
rect 50 143845 62 144821
rect 96 143845 108 144821
rect 50 143833 108 143845
rect -108 143603 -50 143615
rect -108 142627 -96 143603
rect -62 142627 -50 143603
rect -108 142615 -50 142627
rect 50 143603 108 143615
rect 50 142627 62 143603
rect 96 142627 108 143603
rect 50 142615 108 142627
rect -108 142385 -50 142397
rect -108 141409 -96 142385
rect -62 141409 -50 142385
rect -108 141397 -50 141409
rect 50 142385 108 142397
rect 50 141409 62 142385
rect 96 141409 108 142385
rect 50 141397 108 141409
rect -108 141167 -50 141179
rect -108 140191 -96 141167
rect -62 140191 -50 141167
rect -108 140179 -50 140191
rect 50 141167 108 141179
rect 50 140191 62 141167
rect 96 140191 108 141167
rect 50 140179 108 140191
rect -108 139949 -50 139961
rect -108 138973 -96 139949
rect -62 138973 -50 139949
rect -108 138961 -50 138973
rect 50 139949 108 139961
rect 50 138973 62 139949
rect 96 138973 108 139949
rect 50 138961 108 138973
rect -108 138731 -50 138743
rect -108 137755 -96 138731
rect -62 137755 -50 138731
rect -108 137743 -50 137755
rect 50 138731 108 138743
rect 50 137755 62 138731
rect 96 137755 108 138731
rect 50 137743 108 137755
rect -108 137513 -50 137525
rect -108 136537 -96 137513
rect -62 136537 -50 137513
rect -108 136525 -50 136537
rect 50 137513 108 137525
rect 50 136537 62 137513
rect 96 136537 108 137513
rect 50 136525 108 136537
rect -108 136295 -50 136307
rect -108 135319 -96 136295
rect -62 135319 -50 136295
rect -108 135307 -50 135319
rect 50 136295 108 136307
rect 50 135319 62 136295
rect 96 135319 108 136295
rect 50 135307 108 135319
rect -108 135077 -50 135089
rect -108 134101 -96 135077
rect -62 134101 -50 135077
rect -108 134089 -50 134101
rect 50 135077 108 135089
rect 50 134101 62 135077
rect 96 134101 108 135077
rect 50 134089 108 134101
rect -108 133859 -50 133871
rect -108 132883 -96 133859
rect -62 132883 -50 133859
rect -108 132871 -50 132883
rect 50 133859 108 133871
rect 50 132883 62 133859
rect 96 132883 108 133859
rect 50 132871 108 132883
rect -108 132641 -50 132653
rect -108 131665 -96 132641
rect -62 131665 -50 132641
rect -108 131653 -50 131665
rect 50 132641 108 132653
rect 50 131665 62 132641
rect 96 131665 108 132641
rect 50 131653 108 131665
rect -108 131423 -50 131435
rect -108 130447 -96 131423
rect -62 130447 -50 131423
rect -108 130435 -50 130447
rect 50 131423 108 131435
rect 50 130447 62 131423
rect 96 130447 108 131423
rect 50 130435 108 130447
rect -108 130205 -50 130217
rect -108 129229 -96 130205
rect -62 129229 -50 130205
rect -108 129217 -50 129229
rect 50 130205 108 130217
rect 50 129229 62 130205
rect 96 129229 108 130205
rect 50 129217 108 129229
rect -108 128987 -50 128999
rect -108 128011 -96 128987
rect -62 128011 -50 128987
rect -108 127999 -50 128011
rect 50 128987 108 128999
rect 50 128011 62 128987
rect 96 128011 108 128987
rect 50 127999 108 128011
rect -108 127769 -50 127781
rect -108 126793 -96 127769
rect -62 126793 -50 127769
rect -108 126781 -50 126793
rect 50 127769 108 127781
rect 50 126793 62 127769
rect 96 126793 108 127769
rect 50 126781 108 126793
rect -108 126551 -50 126563
rect -108 125575 -96 126551
rect -62 125575 -50 126551
rect -108 125563 -50 125575
rect 50 126551 108 126563
rect 50 125575 62 126551
rect 96 125575 108 126551
rect 50 125563 108 125575
rect -108 125333 -50 125345
rect -108 124357 -96 125333
rect -62 124357 -50 125333
rect -108 124345 -50 124357
rect 50 125333 108 125345
rect 50 124357 62 125333
rect 96 124357 108 125333
rect 50 124345 108 124357
rect -108 124115 -50 124127
rect -108 123139 -96 124115
rect -62 123139 -50 124115
rect -108 123127 -50 123139
rect 50 124115 108 124127
rect 50 123139 62 124115
rect 96 123139 108 124115
rect 50 123127 108 123139
rect -108 122897 -50 122909
rect -108 121921 -96 122897
rect -62 121921 -50 122897
rect -108 121909 -50 121921
rect 50 122897 108 122909
rect 50 121921 62 122897
rect 96 121921 108 122897
rect 50 121909 108 121921
rect -108 121679 -50 121691
rect -108 120703 -96 121679
rect -62 120703 -50 121679
rect -108 120691 -50 120703
rect 50 121679 108 121691
rect 50 120703 62 121679
rect 96 120703 108 121679
rect 50 120691 108 120703
rect -108 120461 -50 120473
rect -108 119485 -96 120461
rect -62 119485 -50 120461
rect -108 119473 -50 119485
rect 50 120461 108 120473
rect 50 119485 62 120461
rect 96 119485 108 120461
rect 50 119473 108 119485
rect -108 119243 -50 119255
rect -108 118267 -96 119243
rect -62 118267 -50 119243
rect -108 118255 -50 118267
rect 50 119243 108 119255
rect 50 118267 62 119243
rect 96 118267 108 119243
rect 50 118255 108 118267
rect -108 118025 -50 118037
rect -108 117049 -96 118025
rect -62 117049 -50 118025
rect -108 117037 -50 117049
rect 50 118025 108 118037
rect 50 117049 62 118025
rect 96 117049 108 118025
rect 50 117037 108 117049
rect -108 116807 -50 116819
rect -108 115831 -96 116807
rect -62 115831 -50 116807
rect -108 115819 -50 115831
rect 50 116807 108 116819
rect 50 115831 62 116807
rect 96 115831 108 116807
rect 50 115819 108 115831
rect -108 115589 -50 115601
rect -108 114613 -96 115589
rect -62 114613 -50 115589
rect -108 114601 -50 114613
rect 50 115589 108 115601
rect 50 114613 62 115589
rect 96 114613 108 115589
rect 50 114601 108 114613
rect -108 114371 -50 114383
rect -108 113395 -96 114371
rect -62 113395 -50 114371
rect -108 113383 -50 113395
rect 50 114371 108 114383
rect 50 113395 62 114371
rect 96 113395 108 114371
rect 50 113383 108 113395
rect -108 113153 -50 113165
rect -108 112177 -96 113153
rect -62 112177 -50 113153
rect -108 112165 -50 112177
rect 50 113153 108 113165
rect 50 112177 62 113153
rect 96 112177 108 113153
rect 50 112165 108 112177
rect -108 111935 -50 111947
rect -108 110959 -96 111935
rect -62 110959 -50 111935
rect -108 110947 -50 110959
rect 50 111935 108 111947
rect 50 110959 62 111935
rect 96 110959 108 111935
rect 50 110947 108 110959
rect -108 110717 -50 110729
rect -108 109741 -96 110717
rect -62 109741 -50 110717
rect -108 109729 -50 109741
rect 50 110717 108 110729
rect 50 109741 62 110717
rect 96 109741 108 110717
rect 50 109729 108 109741
rect -108 109499 -50 109511
rect -108 108523 -96 109499
rect -62 108523 -50 109499
rect -108 108511 -50 108523
rect 50 109499 108 109511
rect 50 108523 62 109499
rect 96 108523 108 109499
rect 50 108511 108 108523
rect -108 108281 -50 108293
rect -108 107305 -96 108281
rect -62 107305 -50 108281
rect -108 107293 -50 107305
rect 50 108281 108 108293
rect 50 107305 62 108281
rect 96 107305 108 108281
rect 50 107293 108 107305
rect -108 107063 -50 107075
rect -108 106087 -96 107063
rect -62 106087 -50 107063
rect -108 106075 -50 106087
rect 50 107063 108 107075
rect 50 106087 62 107063
rect 96 106087 108 107063
rect 50 106075 108 106087
rect -108 105845 -50 105857
rect -108 104869 -96 105845
rect -62 104869 -50 105845
rect -108 104857 -50 104869
rect 50 105845 108 105857
rect 50 104869 62 105845
rect 96 104869 108 105845
rect 50 104857 108 104869
rect -108 104627 -50 104639
rect -108 103651 -96 104627
rect -62 103651 -50 104627
rect -108 103639 -50 103651
rect 50 104627 108 104639
rect 50 103651 62 104627
rect 96 103651 108 104627
rect 50 103639 108 103651
rect -108 103409 -50 103421
rect -108 102433 -96 103409
rect -62 102433 -50 103409
rect -108 102421 -50 102433
rect 50 103409 108 103421
rect 50 102433 62 103409
rect 96 102433 108 103409
rect 50 102421 108 102433
rect -108 102191 -50 102203
rect -108 101215 -96 102191
rect -62 101215 -50 102191
rect -108 101203 -50 101215
rect 50 102191 108 102203
rect 50 101215 62 102191
rect 96 101215 108 102191
rect 50 101203 108 101215
rect -108 100973 -50 100985
rect -108 99997 -96 100973
rect -62 99997 -50 100973
rect -108 99985 -50 99997
rect 50 100973 108 100985
rect 50 99997 62 100973
rect 96 99997 108 100973
rect 50 99985 108 99997
rect -108 99755 -50 99767
rect -108 98779 -96 99755
rect -62 98779 -50 99755
rect -108 98767 -50 98779
rect 50 99755 108 99767
rect 50 98779 62 99755
rect 96 98779 108 99755
rect 50 98767 108 98779
rect -108 98537 -50 98549
rect -108 97561 -96 98537
rect -62 97561 -50 98537
rect -108 97549 -50 97561
rect 50 98537 108 98549
rect 50 97561 62 98537
rect 96 97561 108 98537
rect 50 97549 108 97561
rect -108 97319 -50 97331
rect -108 96343 -96 97319
rect -62 96343 -50 97319
rect -108 96331 -50 96343
rect 50 97319 108 97331
rect 50 96343 62 97319
rect 96 96343 108 97319
rect 50 96331 108 96343
rect -108 96101 -50 96113
rect -108 95125 -96 96101
rect -62 95125 -50 96101
rect -108 95113 -50 95125
rect 50 96101 108 96113
rect 50 95125 62 96101
rect 96 95125 108 96101
rect 50 95113 108 95125
rect -108 94883 -50 94895
rect -108 93907 -96 94883
rect -62 93907 -50 94883
rect -108 93895 -50 93907
rect 50 94883 108 94895
rect 50 93907 62 94883
rect 96 93907 108 94883
rect 50 93895 108 93907
rect -108 93665 -50 93677
rect -108 92689 -96 93665
rect -62 92689 -50 93665
rect -108 92677 -50 92689
rect 50 93665 108 93677
rect 50 92689 62 93665
rect 96 92689 108 93665
rect 50 92677 108 92689
rect -108 92447 -50 92459
rect -108 91471 -96 92447
rect -62 91471 -50 92447
rect -108 91459 -50 91471
rect 50 92447 108 92459
rect 50 91471 62 92447
rect 96 91471 108 92447
rect 50 91459 108 91471
rect -108 91229 -50 91241
rect -108 90253 -96 91229
rect -62 90253 -50 91229
rect -108 90241 -50 90253
rect 50 91229 108 91241
rect 50 90253 62 91229
rect 96 90253 108 91229
rect 50 90241 108 90253
rect -108 90011 -50 90023
rect -108 89035 -96 90011
rect -62 89035 -50 90011
rect -108 89023 -50 89035
rect 50 90011 108 90023
rect 50 89035 62 90011
rect 96 89035 108 90011
rect 50 89023 108 89035
rect -108 88793 -50 88805
rect -108 87817 -96 88793
rect -62 87817 -50 88793
rect -108 87805 -50 87817
rect 50 88793 108 88805
rect 50 87817 62 88793
rect 96 87817 108 88793
rect 50 87805 108 87817
rect -108 87575 -50 87587
rect -108 86599 -96 87575
rect -62 86599 -50 87575
rect -108 86587 -50 86599
rect 50 87575 108 87587
rect 50 86599 62 87575
rect 96 86599 108 87575
rect 50 86587 108 86599
rect -108 86357 -50 86369
rect -108 85381 -96 86357
rect -62 85381 -50 86357
rect -108 85369 -50 85381
rect 50 86357 108 86369
rect 50 85381 62 86357
rect 96 85381 108 86357
rect 50 85369 108 85381
rect -108 85139 -50 85151
rect -108 84163 -96 85139
rect -62 84163 -50 85139
rect -108 84151 -50 84163
rect 50 85139 108 85151
rect 50 84163 62 85139
rect 96 84163 108 85139
rect 50 84151 108 84163
rect -108 83921 -50 83933
rect -108 82945 -96 83921
rect -62 82945 -50 83921
rect -108 82933 -50 82945
rect 50 83921 108 83933
rect 50 82945 62 83921
rect 96 82945 108 83921
rect 50 82933 108 82945
rect -108 82703 -50 82715
rect -108 81727 -96 82703
rect -62 81727 -50 82703
rect -108 81715 -50 81727
rect 50 82703 108 82715
rect 50 81727 62 82703
rect 96 81727 108 82703
rect 50 81715 108 81727
rect -108 81485 -50 81497
rect -108 80509 -96 81485
rect -62 80509 -50 81485
rect -108 80497 -50 80509
rect 50 81485 108 81497
rect 50 80509 62 81485
rect 96 80509 108 81485
rect 50 80497 108 80509
rect -108 80267 -50 80279
rect -108 79291 -96 80267
rect -62 79291 -50 80267
rect -108 79279 -50 79291
rect 50 80267 108 80279
rect 50 79291 62 80267
rect 96 79291 108 80267
rect 50 79279 108 79291
rect -108 79049 -50 79061
rect -108 78073 -96 79049
rect -62 78073 -50 79049
rect -108 78061 -50 78073
rect 50 79049 108 79061
rect 50 78073 62 79049
rect 96 78073 108 79049
rect 50 78061 108 78073
rect -108 77831 -50 77843
rect -108 76855 -96 77831
rect -62 76855 -50 77831
rect -108 76843 -50 76855
rect 50 77831 108 77843
rect 50 76855 62 77831
rect 96 76855 108 77831
rect 50 76843 108 76855
rect -108 76613 -50 76625
rect -108 75637 -96 76613
rect -62 75637 -50 76613
rect -108 75625 -50 75637
rect 50 76613 108 76625
rect 50 75637 62 76613
rect 96 75637 108 76613
rect 50 75625 108 75637
rect -108 75395 -50 75407
rect -108 74419 -96 75395
rect -62 74419 -50 75395
rect -108 74407 -50 74419
rect 50 75395 108 75407
rect 50 74419 62 75395
rect 96 74419 108 75395
rect 50 74407 108 74419
rect -108 74177 -50 74189
rect -108 73201 -96 74177
rect -62 73201 -50 74177
rect -108 73189 -50 73201
rect 50 74177 108 74189
rect 50 73201 62 74177
rect 96 73201 108 74177
rect 50 73189 108 73201
rect -108 72959 -50 72971
rect -108 71983 -96 72959
rect -62 71983 -50 72959
rect -108 71971 -50 71983
rect 50 72959 108 72971
rect 50 71983 62 72959
rect 96 71983 108 72959
rect 50 71971 108 71983
rect -108 71741 -50 71753
rect -108 70765 -96 71741
rect -62 70765 -50 71741
rect -108 70753 -50 70765
rect 50 71741 108 71753
rect 50 70765 62 71741
rect 96 70765 108 71741
rect 50 70753 108 70765
rect -108 70523 -50 70535
rect -108 69547 -96 70523
rect -62 69547 -50 70523
rect -108 69535 -50 69547
rect 50 70523 108 70535
rect 50 69547 62 70523
rect 96 69547 108 70523
rect 50 69535 108 69547
rect -108 69305 -50 69317
rect -108 68329 -96 69305
rect -62 68329 -50 69305
rect -108 68317 -50 68329
rect 50 69305 108 69317
rect 50 68329 62 69305
rect 96 68329 108 69305
rect 50 68317 108 68329
rect -108 68087 -50 68099
rect -108 67111 -96 68087
rect -62 67111 -50 68087
rect -108 67099 -50 67111
rect 50 68087 108 68099
rect 50 67111 62 68087
rect 96 67111 108 68087
rect 50 67099 108 67111
rect -108 66869 -50 66881
rect -108 65893 -96 66869
rect -62 65893 -50 66869
rect -108 65881 -50 65893
rect 50 66869 108 66881
rect 50 65893 62 66869
rect 96 65893 108 66869
rect 50 65881 108 65893
rect -108 65651 -50 65663
rect -108 64675 -96 65651
rect -62 64675 -50 65651
rect -108 64663 -50 64675
rect 50 65651 108 65663
rect 50 64675 62 65651
rect 96 64675 108 65651
rect 50 64663 108 64675
rect -108 64433 -50 64445
rect -108 63457 -96 64433
rect -62 63457 -50 64433
rect -108 63445 -50 63457
rect 50 64433 108 64445
rect 50 63457 62 64433
rect 96 63457 108 64433
rect 50 63445 108 63457
rect -108 63215 -50 63227
rect -108 62239 -96 63215
rect -62 62239 -50 63215
rect -108 62227 -50 62239
rect 50 63215 108 63227
rect 50 62239 62 63215
rect 96 62239 108 63215
rect 50 62227 108 62239
rect -108 61997 -50 62009
rect -108 61021 -96 61997
rect -62 61021 -50 61997
rect -108 61009 -50 61021
rect 50 61997 108 62009
rect 50 61021 62 61997
rect 96 61021 108 61997
rect 50 61009 108 61021
rect -108 60779 -50 60791
rect -108 59803 -96 60779
rect -62 59803 -50 60779
rect -108 59791 -50 59803
rect 50 60779 108 60791
rect 50 59803 62 60779
rect 96 59803 108 60779
rect 50 59791 108 59803
rect -108 59561 -50 59573
rect -108 58585 -96 59561
rect -62 58585 -50 59561
rect -108 58573 -50 58585
rect 50 59561 108 59573
rect 50 58585 62 59561
rect 96 58585 108 59561
rect 50 58573 108 58585
rect -108 58343 -50 58355
rect -108 57367 -96 58343
rect -62 57367 -50 58343
rect -108 57355 -50 57367
rect 50 58343 108 58355
rect 50 57367 62 58343
rect 96 57367 108 58343
rect 50 57355 108 57367
rect -108 57125 -50 57137
rect -108 56149 -96 57125
rect -62 56149 -50 57125
rect -108 56137 -50 56149
rect 50 57125 108 57137
rect 50 56149 62 57125
rect 96 56149 108 57125
rect 50 56137 108 56149
rect -108 55907 -50 55919
rect -108 54931 -96 55907
rect -62 54931 -50 55907
rect -108 54919 -50 54931
rect 50 55907 108 55919
rect 50 54931 62 55907
rect 96 54931 108 55907
rect 50 54919 108 54931
rect -108 54689 -50 54701
rect -108 53713 -96 54689
rect -62 53713 -50 54689
rect -108 53701 -50 53713
rect 50 54689 108 54701
rect 50 53713 62 54689
rect 96 53713 108 54689
rect 50 53701 108 53713
rect -108 53471 -50 53483
rect -108 52495 -96 53471
rect -62 52495 -50 53471
rect -108 52483 -50 52495
rect 50 53471 108 53483
rect 50 52495 62 53471
rect 96 52495 108 53471
rect 50 52483 108 52495
rect -108 52253 -50 52265
rect -108 51277 -96 52253
rect -62 51277 -50 52253
rect -108 51265 -50 51277
rect 50 52253 108 52265
rect 50 51277 62 52253
rect 96 51277 108 52253
rect 50 51265 108 51277
rect -108 51035 -50 51047
rect -108 50059 -96 51035
rect -62 50059 -50 51035
rect -108 50047 -50 50059
rect 50 51035 108 51047
rect 50 50059 62 51035
rect 96 50059 108 51035
rect 50 50047 108 50059
rect -108 49817 -50 49829
rect -108 48841 -96 49817
rect -62 48841 -50 49817
rect -108 48829 -50 48841
rect 50 49817 108 49829
rect 50 48841 62 49817
rect 96 48841 108 49817
rect 50 48829 108 48841
rect -108 48599 -50 48611
rect -108 47623 -96 48599
rect -62 47623 -50 48599
rect -108 47611 -50 47623
rect 50 48599 108 48611
rect 50 47623 62 48599
rect 96 47623 108 48599
rect 50 47611 108 47623
rect -108 47381 -50 47393
rect -108 46405 -96 47381
rect -62 46405 -50 47381
rect -108 46393 -50 46405
rect 50 47381 108 47393
rect 50 46405 62 47381
rect 96 46405 108 47381
rect 50 46393 108 46405
rect -108 46163 -50 46175
rect -108 45187 -96 46163
rect -62 45187 -50 46163
rect -108 45175 -50 45187
rect 50 46163 108 46175
rect 50 45187 62 46163
rect 96 45187 108 46163
rect 50 45175 108 45187
rect -108 44945 -50 44957
rect -108 43969 -96 44945
rect -62 43969 -50 44945
rect -108 43957 -50 43969
rect 50 44945 108 44957
rect 50 43969 62 44945
rect 96 43969 108 44945
rect 50 43957 108 43969
rect -108 43727 -50 43739
rect -108 42751 -96 43727
rect -62 42751 -50 43727
rect -108 42739 -50 42751
rect 50 43727 108 43739
rect 50 42751 62 43727
rect 96 42751 108 43727
rect 50 42739 108 42751
rect -108 42509 -50 42521
rect -108 41533 -96 42509
rect -62 41533 -50 42509
rect -108 41521 -50 41533
rect 50 42509 108 42521
rect 50 41533 62 42509
rect 96 41533 108 42509
rect 50 41521 108 41533
rect -108 41291 -50 41303
rect -108 40315 -96 41291
rect -62 40315 -50 41291
rect -108 40303 -50 40315
rect 50 41291 108 41303
rect 50 40315 62 41291
rect 96 40315 108 41291
rect 50 40303 108 40315
rect -108 40073 -50 40085
rect -108 39097 -96 40073
rect -62 39097 -50 40073
rect -108 39085 -50 39097
rect 50 40073 108 40085
rect 50 39097 62 40073
rect 96 39097 108 40073
rect 50 39085 108 39097
rect -108 38855 -50 38867
rect -108 37879 -96 38855
rect -62 37879 -50 38855
rect -108 37867 -50 37879
rect 50 38855 108 38867
rect 50 37879 62 38855
rect 96 37879 108 38855
rect 50 37867 108 37879
rect -108 37637 -50 37649
rect -108 36661 -96 37637
rect -62 36661 -50 37637
rect -108 36649 -50 36661
rect 50 37637 108 37649
rect 50 36661 62 37637
rect 96 36661 108 37637
rect 50 36649 108 36661
rect -108 36419 -50 36431
rect -108 35443 -96 36419
rect -62 35443 -50 36419
rect -108 35431 -50 35443
rect 50 36419 108 36431
rect 50 35443 62 36419
rect 96 35443 108 36419
rect 50 35431 108 35443
rect -108 35201 -50 35213
rect -108 34225 -96 35201
rect -62 34225 -50 35201
rect -108 34213 -50 34225
rect 50 35201 108 35213
rect 50 34225 62 35201
rect 96 34225 108 35201
rect 50 34213 108 34225
rect -108 33983 -50 33995
rect -108 33007 -96 33983
rect -62 33007 -50 33983
rect -108 32995 -50 33007
rect 50 33983 108 33995
rect 50 33007 62 33983
rect 96 33007 108 33983
rect 50 32995 108 33007
rect -108 32765 -50 32777
rect -108 31789 -96 32765
rect -62 31789 -50 32765
rect -108 31777 -50 31789
rect 50 32765 108 32777
rect 50 31789 62 32765
rect 96 31789 108 32765
rect 50 31777 108 31789
rect -108 31547 -50 31559
rect -108 30571 -96 31547
rect -62 30571 -50 31547
rect -108 30559 -50 30571
rect 50 31547 108 31559
rect 50 30571 62 31547
rect 96 30571 108 31547
rect 50 30559 108 30571
rect -108 30329 -50 30341
rect -108 29353 -96 30329
rect -62 29353 -50 30329
rect -108 29341 -50 29353
rect 50 30329 108 30341
rect 50 29353 62 30329
rect 96 29353 108 30329
rect 50 29341 108 29353
rect -108 29111 -50 29123
rect -108 28135 -96 29111
rect -62 28135 -50 29111
rect -108 28123 -50 28135
rect 50 29111 108 29123
rect 50 28135 62 29111
rect 96 28135 108 29111
rect 50 28123 108 28135
rect -108 27893 -50 27905
rect -108 26917 -96 27893
rect -62 26917 -50 27893
rect -108 26905 -50 26917
rect 50 27893 108 27905
rect 50 26917 62 27893
rect 96 26917 108 27893
rect 50 26905 108 26917
rect -108 26675 -50 26687
rect -108 25699 -96 26675
rect -62 25699 -50 26675
rect -108 25687 -50 25699
rect 50 26675 108 26687
rect 50 25699 62 26675
rect 96 25699 108 26675
rect 50 25687 108 25699
rect -108 25457 -50 25469
rect -108 24481 -96 25457
rect -62 24481 -50 25457
rect -108 24469 -50 24481
rect 50 25457 108 25469
rect 50 24481 62 25457
rect 96 24481 108 25457
rect 50 24469 108 24481
rect -108 24239 -50 24251
rect -108 23263 -96 24239
rect -62 23263 -50 24239
rect -108 23251 -50 23263
rect 50 24239 108 24251
rect 50 23263 62 24239
rect 96 23263 108 24239
rect 50 23251 108 23263
rect -108 23021 -50 23033
rect -108 22045 -96 23021
rect -62 22045 -50 23021
rect -108 22033 -50 22045
rect 50 23021 108 23033
rect 50 22045 62 23021
rect 96 22045 108 23021
rect 50 22033 108 22045
rect -108 21803 -50 21815
rect -108 20827 -96 21803
rect -62 20827 -50 21803
rect -108 20815 -50 20827
rect 50 21803 108 21815
rect 50 20827 62 21803
rect 96 20827 108 21803
rect 50 20815 108 20827
rect -108 20585 -50 20597
rect -108 19609 -96 20585
rect -62 19609 -50 20585
rect -108 19597 -50 19609
rect 50 20585 108 20597
rect 50 19609 62 20585
rect 96 19609 108 20585
rect 50 19597 108 19609
rect -108 19367 -50 19379
rect -108 18391 -96 19367
rect -62 18391 -50 19367
rect -108 18379 -50 18391
rect 50 19367 108 19379
rect 50 18391 62 19367
rect 96 18391 108 19367
rect 50 18379 108 18391
rect -108 18149 -50 18161
rect -108 17173 -96 18149
rect -62 17173 -50 18149
rect -108 17161 -50 17173
rect 50 18149 108 18161
rect 50 17173 62 18149
rect 96 17173 108 18149
rect 50 17161 108 17173
rect -108 16931 -50 16943
rect -108 15955 -96 16931
rect -62 15955 -50 16931
rect -108 15943 -50 15955
rect 50 16931 108 16943
rect 50 15955 62 16931
rect 96 15955 108 16931
rect 50 15943 108 15955
rect -108 15713 -50 15725
rect -108 14737 -96 15713
rect -62 14737 -50 15713
rect -108 14725 -50 14737
rect 50 15713 108 15725
rect 50 14737 62 15713
rect 96 14737 108 15713
rect 50 14725 108 14737
rect -108 14495 -50 14507
rect -108 13519 -96 14495
rect -62 13519 -50 14495
rect -108 13507 -50 13519
rect 50 14495 108 14507
rect 50 13519 62 14495
rect 96 13519 108 14495
rect 50 13507 108 13519
rect -108 13277 -50 13289
rect -108 12301 -96 13277
rect -62 12301 -50 13277
rect -108 12289 -50 12301
rect 50 13277 108 13289
rect 50 12301 62 13277
rect 96 12301 108 13277
rect 50 12289 108 12301
rect -108 12059 -50 12071
rect -108 11083 -96 12059
rect -62 11083 -50 12059
rect -108 11071 -50 11083
rect 50 12059 108 12071
rect 50 11083 62 12059
rect 96 11083 108 12059
rect 50 11071 108 11083
rect -108 10841 -50 10853
rect -108 9865 -96 10841
rect -62 9865 -50 10841
rect -108 9853 -50 9865
rect 50 10841 108 10853
rect 50 9865 62 10841
rect 96 9865 108 10841
rect 50 9853 108 9865
rect -108 9623 -50 9635
rect -108 8647 -96 9623
rect -62 8647 -50 9623
rect -108 8635 -50 8647
rect 50 9623 108 9635
rect 50 8647 62 9623
rect 96 8647 108 9623
rect 50 8635 108 8647
rect -108 8405 -50 8417
rect -108 7429 -96 8405
rect -62 7429 -50 8405
rect -108 7417 -50 7429
rect 50 8405 108 8417
rect 50 7429 62 8405
rect 96 7429 108 8405
rect 50 7417 108 7429
rect -108 7187 -50 7199
rect -108 6211 -96 7187
rect -62 6211 -50 7187
rect -108 6199 -50 6211
rect 50 7187 108 7199
rect 50 6211 62 7187
rect 96 6211 108 7187
rect 50 6199 108 6211
rect -108 5969 -50 5981
rect -108 4993 -96 5969
rect -62 4993 -50 5969
rect -108 4981 -50 4993
rect 50 5969 108 5981
rect 50 4993 62 5969
rect 96 4993 108 5969
rect 50 4981 108 4993
rect -108 4751 -50 4763
rect -108 3775 -96 4751
rect -62 3775 -50 4751
rect -108 3763 -50 3775
rect 50 4751 108 4763
rect 50 3775 62 4751
rect 96 3775 108 4751
rect 50 3763 108 3775
rect -108 3533 -50 3545
rect -108 2557 -96 3533
rect -62 2557 -50 3533
rect -108 2545 -50 2557
rect 50 3533 108 3545
rect 50 2557 62 3533
rect 96 2557 108 3533
rect 50 2545 108 2557
rect -108 2315 -50 2327
rect -108 1339 -96 2315
rect -62 1339 -50 2315
rect -108 1327 -50 1339
rect 50 2315 108 2327
rect 50 1339 62 2315
rect 96 1339 108 2315
rect 50 1327 108 1339
rect -108 1097 -50 1109
rect -108 121 -96 1097
rect -62 121 -50 1097
rect -108 109 -50 121
rect 50 1097 108 1109
rect 50 121 62 1097
rect 96 121 108 1097
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -1097 -96 -121
rect -62 -1097 -50 -121
rect -108 -1109 -50 -1097
rect 50 -121 108 -109
rect 50 -1097 62 -121
rect 96 -1097 108 -121
rect 50 -1109 108 -1097
rect -108 -1339 -50 -1327
rect -108 -2315 -96 -1339
rect -62 -2315 -50 -1339
rect -108 -2327 -50 -2315
rect 50 -1339 108 -1327
rect 50 -2315 62 -1339
rect 96 -2315 108 -1339
rect 50 -2327 108 -2315
rect -108 -2557 -50 -2545
rect -108 -3533 -96 -2557
rect -62 -3533 -50 -2557
rect -108 -3545 -50 -3533
rect 50 -2557 108 -2545
rect 50 -3533 62 -2557
rect 96 -3533 108 -2557
rect 50 -3545 108 -3533
rect -108 -3775 -50 -3763
rect -108 -4751 -96 -3775
rect -62 -4751 -50 -3775
rect -108 -4763 -50 -4751
rect 50 -3775 108 -3763
rect 50 -4751 62 -3775
rect 96 -4751 108 -3775
rect 50 -4763 108 -4751
rect -108 -4993 -50 -4981
rect -108 -5969 -96 -4993
rect -62 -5969 -50 -4993
rect -108 -5981 -50 -5969
rect 50 -4993 108 -4981
rect 50 -5969 62 -4993
rect 96 -5969 108 -4993
rect 50 -5981 108 -5969
rect -108 -6211 -50 -6199
rect -108 -7187 -96 -6211
rect -62 -7187 -50 -6211
rect -108 -7199 -50 -7187
rect 50 -6211 108 -6199
rect 50 -7187 62 -6211
rect 96 -7187 108 -6211
rect 50 -7199 108 -7187
rect -108 -7429 -50 -7417
rect -108 -8405 -96 -7429
rect -62 -8405 -50 -7429
rect -108 -8417 -50 -8405
rect 50 -7429 108 -7417
rect 50 -8405 62 -7429
rect 96 -8405 108 -7429
rect 50 -8417 108 -8405
rect -108 -8647 -50 -8635
rect -108 -9623 -96 -8647
rect -62 -9623 -50 -8647
rect -108 -9635 -50 -9623
rect 50 -8647 108 -8635
rect 50 -9623 62 -8647
rect 96 -9623 108 -8647
rect 50 -9635 108 -9623
rect -108 -9865 -50 -9853
rect -108 -10841 -96 -9865
rect -62 -10841 -50 -9865
rect -108 -10853 -50 -10841
rect 50 -9865 108 -9853
rect 50 -10841 62 -9865
rect 96 -10841 108 -9865
rect 50 -10853 108 -10841
rect -108 -11083 -50 -11071
rect -108 -12059 -96 -11083
rect -62 -12059 -50 -11083
rect -108 -12071 -50 -12059
rect 50 -11083 108 -11071
rect 50 -12059 62 -11083
rect 96 -12059 108 -11083
rect 50 -12071 108 -12059
rect -108 -12301 -50 -12289
rect -108 -13277 -96 -12301
rect -62 -13277 -50 -12301
rect -108 -13289 -50 -13277
rect 50 -12301 108 -12289
rect 50 -13277 62 -12301
rect 96 -13277 108 -12301
rect 50 -13289 108 -13277
rect -108 -13519 -50 -13507
rect -108 -14495 -96 -13519
rect -62 -14495 -50 -13519
rect -108 -14507 -50 -14495
rect 50 -13519 108 -13507
rect 50 -14495 62 -13519
rect 96 -14495 108 -13519
rect 50 -14507 108 -14495
rect -108 -14737 -50 -14725
rect -108 -15713 -96 -14737
rect -62 -15713 -50 -14737
rect -108 -15725 -50 -15713
rect 50 -14737 108 -14725
rect 50 -15713 62 -14737
rect 96 -15713 108 -14737
rect 50 -15725 108 -15713
rect -108 -15955 -50 -15943
rect -108 -16931 -96 -15955
rect -62 -16931 -50 -15955
rect -108 -16943 -50 -16931
rect 50 -15955 108 -15943
rect 50 -16931 62 -15955
rect 96 -16931 108 -15955
rect 50 -16943 108 -16931
rect -108 -17173 -50 -17161
rect -108 -18149 -96 -17173
rect -62 -18149 -50 -17173
rect -108 -18161 -50 -18149
rect 50 -17173 108 -17161
rect 50 -18149 62 -17173
rect 96 -18149 108 -17173
rect 50 -18161 108 -18149
rect -108 -18391 -50 -18379
rect -108 -19367 -96 -18391
rect -62 -19367 -50 -18391
rect -108 -19379 -50 -19367
rect 50 -18391 108 -18379
rect 50 -19367 62 -18391
rect 96 -19367 108 -18391
rect 50 -19379 108 -19367
rect -108 -19609 -50 -19597
rect -108 -20585 -96 -19609
rect -62 -20585 -50 -19609
rect -108 -20597 -50 -20585
rect 50 -19609 108 -19597
rect 50 -20585 62 -19609
rect 96 -20585 108 -19609
rect 50 -20597 108 -20585
rect -108 -20827 -50 -20815
rect -108 -21803 -96 -20827
rect -62 -21803 -50 -20827
rect -108 -21815 -50 -21803
rect 50 -20827 108 -20815
rect 50 -21803 62 -20827
rect 96 -21803 108 -20827
rect 50 -21815 108 -21803
rect -108 -22045 -50 -22033
rect -108 -23021 -96 -22045
rect -62 -23021 -50 -22045
rect -108 -23033 -50 -23021
rect 50 -22045 108 -22033
rect 50 -23021 62 -22045
rect 96 -23021 108 -22045
rect 50 -23033 108 -23021
rect -108 -23263 -50 -23251
rect -108 -24239 -96 -23263
rect -62 -24239 -50 -23263
rect -108 -24251 -50 -24239
rect 50 -23263 108 -23251
rect 50 -24239 62 -23263
rect 96 -24239 108 -23263
rect 50 -24251 108 -24239
rect -108 -24481 -50 -24469
rect -108 -25457 -96 -24481
rect -62 -25457 -50 -24481
rect -108 -25469 -50 -25457
rect 50 -24481 108 -24469
rect 50 -25457 62 -24481
rect 96 -25457 108 -24481
rect 50 -25469 108 -25457
rect -108 -25699 -50 -25687
rect -108 -26675 -96 -25699
rect -62 -26675 -50 -25699
rect -108 -26687 -50 -26675
rect 50 -25699 108 -25687
rect 50 -26675 62 -25699
rect 96 -26675 108 -25699
rect 50 -26687 108 -26675
rect -108 -26917 -50 -26905
rect -108 -27893 -96 -26917
rect -62 -27893 -50 -26917
rect -108 -27905 -50 -27893
rect 50 -26917 108 -26905
rect 50 -27893 62 -26917
rect 96 -27893 108 -26917
rect 50 -27905 108 -27893
rect -108 -28135 -50 -28123
rect -108 -29111 -96 -28135
rect -62 -29111 -50 -28135
rect -108 -29123 -50 -29111
rect 50 -28135 108 -28123
rect 50 -29111 62 -28135
rect 96 -29111 108 -28135
rect 50 -29123 108 -29111
rect -108 -29353 -50 -29341
rect -108 -30329 -96 -29353
rect -62 -30329 -50 -29353
rect -108 -30341 -50 -30329
rect 50 -29353 108 -29341
rect 50 -30329 62 -29353
rect 96 -30329 108 -29353
rect 50 -30341 108 -30329
rect -108 -30571 -50 -30559
rect -108 -31547 -96 -30571
rect -62 -31547 -50 -30571
rect -108 -31559 -50 -31547
rect 50 -30571 108 -30559
rect 50 -31547 62 -30571
rect 96 -31547 108 -30571
rect 50 -31559 108 -31547
rect -108 -31789 -50 -31777
rect -108 -32765 -96 -31789
rect -62 -32765 -50 -31789
rect -108 -32777 -50 -32765
rect 50 -31789 108 -31777
rect 50 -32765 62 -31789
rect 96 -32765 108 -31789
rect 50 -32777 108 -32765
rect -108 -33007 -50 -32995
rect -108 -33983 -96 -33007
rect -62 -33983 -50 -33007
rect -108 -33995 -50 -33983
rect 50 -33007 108 -32995
rect 50 -33983 62 -33007
rect 96 -33983 108 -33007
rect 50 -33995 108 -33983
rect -108 -34225 -50 -34213
rect -108 -35201 -96 -34225
rect -62 -35201 -50 -34225
rect -108 -35213 -50 -35201
rect 50 -34225 108 -34213
rect 50 -35201 62 -34225
rect 96 -35201 108 -34225
rect 50 -35213 108 -35201
rect -108 -35443 -50 -35431
rect -108 -36419 -96 -35443
rect -62 -36419 -50 -35443
rect -108 -36431 -50 -36419
rect 50 -35443 108 -35431
rect 50 -36419 62 -35443
rect 96 -36419 108 -35443
rect 50 -36431 108 -36419
rect -108 -36661 -50 -36649
rect -108 -37637 -96 -36661
rect -62 -37637 -50 -36661
rect -108 -37649 -50 -37637
rect 50 -36661 108 -36649
rect 50 -37637 62 -36661
rect 96 -37637 108 -36661
rect 50 -37649 108 -37637
rect -108 -37879 -50 -37867
rect -108 -38855 -96 -37879
rect -62 -38855 -50 -37879
rect -108 -38867 -50 -38855
rect 50 -37879 108 -37867
rect 50 -38855 62 -37879
rect 96 -38855 108 -37879
rect 50 -38867 108 -38855
rect -108 -39097 -50 -39085
rect -108 -40073 -96 -39097
rect -62 -40073 -50 -39097
rect -108 -40085 -50 -40073
rect 50 -39097 108 -39085
rect 50 -40073 62 -39097
rect 96 -40073 108 -39097
rect 50 -40085 108 -40073
rect -108 -40315 -50 -40303
rect -108 -41291 -96 -40315
rect -62 -41291 -50 -40315
rect -108 -41303 -50 -41291
rect 50 -40315 108 -40303
rect 50 -41291 62 -40315
rect 96 -41291 108 -40315
rect 50 -41303 108 -41291
rect -108 -41533 -50 -41521
rect -108 -42509 -96 -41533
rect -62 -42509 -50 -41533
rect -108 -42521 -50 -42509
rect 50 -41533 108 -41521
rect 50 -42509 62 -41533
rect 96 -42509 108 -41533
rect 50 -42521 108 -42509
rect -108 -42751 -50 -42739
rect -108 -43727 -96 -42751
rect -62 -43727 -50 -42751
rect -108 -43739 -50 -43727
rect 50 -42751 108 -42739
rect 50 -43727 62 -42751
rect 96 -43727 108 -42751
rect 50 -43739 108 -43727
rect -108 -43969 -50 -43957
rect -108 -44945 -96 -43969
rect -62 -44945 -50 -43969
rect -108 -44957 -50 -44945
rect 50 -43969 108 -43957
rect 50 -44945 62 -43969
rect 96 -44945 108 -43969
rect 50 -44957 108 -44945
rect -108 -45187 -50 -45175
rect -108 -46163 -96 -45187
rect -62 -46163 -50 -45187
rect -108 -46175 -50 -46163
rect 50 -45187 108 -45175
rect 50 -46163 62 -45187
rect 96 -46163 108 -45187
rect 50 -46175 108 -46163
rect -108 -46405 -50 -46393
rect -108 -47381 -96 -46405
rect -62 -47381 -50 -46405
rect -108 -47393 -50 -47381
rect 50 -46405 108 -46393
rect 50 -47381 62 -46405
rect 96 -47381 108 -46405
rect 50 -47393 108 -47381
rect -108 -47623 -50 -47611
rect -108 -48599 -96 -47623
rect -62 -48599 -50 -47623
rect -108 -48611 -50 -48599
rect 50 -47623 108 -47611
rect 50 -48599 62 -47623
rect 96 -48599 108 -47623
rect 50 -48611 108 -48599
rect -108 -48841 -50 -48829
rect -108 -49817 -96 -48841
rect -62 -49817 -50 -48841
rect -108 -49829 -50 -49817
rect 50 -48841 108 -48829
rect 50 -49817 62 -48841
rect 96 -49817 108 -48841
rect 50 -49829 108 -49817
rect -108 -50059 -50 -50047
rect -108 -51035 -96 -50059
rect -62 -51035 -50 -50059
rect -108 -51047 -50 -51035
rect 50 -50059 108 -50047
rect 50 -51035 62 -50059
rect 96 -51035 108 -50059
rect 50 -51047 108 -51035
rect -108 -51277 -50 -51265
rect -108 -52253 -96 -51277
rect -62 -52253 -50 -51277
rect -108 -52265 -50 -52253
rect 50 -51277 108 -51265
rect 50 -52253 62 -51277
rect 96 -52253 108 -51277
rect 50 -52265 108 -52253
rect -108 -52495 -50 -52483
rect -108 -53471 -96 -52495
rect -62 -53471 -50 -52495
rect -108 -53483 -50 -53471
rect 50 -52495 108 -52483
rect 50 -53471 62 -52495
rect 96 -53471 108 -52495
rect 50 -53483 108 -53471
rect -108 -53713 -50 -53701
rect -108 -54689 -96 -53713
rect -62 -54689 -50 -53713
rect -108 -54701 -50 -54689
rect 50 -53713 108 -53701
rect 50 -54689 62 -53713
rect 96 -54689 108 -53713
rect 50 -54701 108 -54689
rect -108 -54931 -50 -54919
rect -108 -55907 -96 -54931
rect -62 -55907 -50 -54931
rect -108 -55919 -50 -55907
rect 50 -54931 108 -54919
rect 50 -55907 62 -54931
rect 96 -55907 108 -54931
rect 50 -55919 108 -55907
rect -108 -56149 -50 -56137
rect -108 -57125 -96 -56149
rect -62 -57125 -50 -56149
rect -108 -57137 -50 -57125
rect 50 -56149 108 -56137
rect 50 -57125 62 -56149
rect 96 -57125 108 -56149
rect 50 -57137 108 -57125
rect -108 -57367 -50 -57355
rect -108 -58343 -96 -57367
rect -62 -58343 -50 -57367
rect -108 -58355 -50 -58343
rect 50 -57367 108 -57355
rect 50 -58343 62 -57367
rect 96 -58343 108 -57367
rect 50 -58355 108 -58343
rect -108 -58585 -50 -58573
rect -108 -59561 -96 -58585
rect -62 -59561 -50 -58585
rect -108 -59573 -50 -59561
rect 50 -58585 108 -58573
rect 50 -59561 62 -58585
rect 96 -59561 108 -58585
rect 50 -59573 108 -59561
rect -108 -59803 -50 -59791
rect -108 -60779 -96 -59803
rect -62 -60779 -50 -59803
rect -108 -60791 -50 -60779
rect 50 -59803 108 -59791
rect 50 -60779 62 -59803
rect 96 -60779 108 -59803
rect 50 -60791 108 -60779
rect -108 -61021 -50 -61009
rect -108 -61997 -96 -61021
rect -62 -61997 -50 -61021
rect -108 -62009 -50 -61997
rect 50 -61021 108 -61009
rect 50 -61997 62 -61021
rect 96 -61997 108 -61021
rect 50 -62009 108 -61997
rect -108 -62239 -50 -62227
rect -108 -63215 -96 -62239
rect -62 -63215 -50 -62239
rect -108 -63227 -50 -63215
rect 50 -62239 108 -62227
rect 50 -63215 62 -62239
rect 96 -63215 108 -62239
rect 50 -63227 108 -63215
rect -108 -63457 -50 -63445
rect -108 -64433 -96 -63457
rect -62 -64433 -50 -63457
rect -108 -64445 -50 -64433
rect 50 -63457 108 -63445
rect 50 -64433 62 -63457
rect 96 -64433 108 -63457
rect 50 -64445 108 -64433
rect -108 -64675 -50 -64663
rect -108 -65651 -96 -64675
rect -62 -65651 -50 -64675
rect -108 -65663 -50 -65651
rect 50 -64675 108 -64663
rect 50 -65651 62 -64675
rect 96 -65651 108 -64675
rect 50 -65663 108 -65651
rect -108 -65893 -50 -65881
rect -108 -66869 -96 -65893
rect -62 -66869 -50 -65893
rect -108 -66881 -50 -66869
rect 50 -65893 108 -65881
rect 50 -66869 62 -65893
rect 96 -66869 108 -65893
rect 50 -66881 108 -66869
rect -108 -67111 -50 -67099
rect -108 -68087 -96 -67111
rect -62 -68087 -50 -67111
rect -108 -68099 -50 -68087
rect 50 -67111 108 -67099
rect 50 -68087 62 -67111
rect 96 -68087 108 -67111
rect 50 -68099 108 -68087
rect -108 -68329 -50 -68317
rect -108 -69305 -96 -68329
rect -62 -69305 -50 -68329
rect -108 -69317 -50 -69305
rect 50 -68329 108 -68317
rect 50 -69305 62 -68329
rect 96 -69305 108 -68329
rect 50 -69317 108 -69305
rect -108 -69547 -50 -69535
rect -108 -70523 -96 -69547
rect -62 -70523 -50 -69547
rect -108 -70535 -50 -70523
rect 50 -69547 108 -69535
rect 50 -70523 62 -69547
rect 96 -70523 108 -69547
rect 50 -70535 108 -70523
rect -108 -70765 -50 -70753
rect -108 -71741 -96 -70765
rect -62 -71741 -50 -70765
rect -108 -71753 -50 -71741
rect 50 -70765 108 -70753
rect 50 -71741 62 -70765
rect 96 -71741 108 -70765
rect 50 -71753 108 -71741
rect -108 -71983 -50 -71971
rect -108 -72959 -96 -71983
rect -62 -72959 -50 -71983
rect -108 -72971 -50 -72959
rect 50 -71983 108 -71971
rect 50 -72959 62 -71983
rect 96 -72959 108 -71983
rect 50 -72971 108 -72959
rect -108 -73201 -50 -73189
rect -108 -74177 -96 -73201
rect -62 -74177 -50 -73201
rect -108 -74189 -50 -74177
rect 50 -73201 108 -73189
rect 50 -74177 62 -73201
rect 96 -74177 108 -73201
rect 50 -74189 108 -74177
rect -108 -74419 -50 -74407
rect -108 -75395 -96 -74419
rect -62 -75395 -50 -74419
rect -108 -75407 -50 -75395
rect 50 -74419 108 -74407
rect 50 -75395 62 -74419
rect 96 -75395 108 -74419
rect 50 -75407 108 -75395
rect -108 -75637 -50 -75625
rect -108 -76613 -96 -75637
rect -62 -76613 -50 -75637
rect -108 -76625 -50 -76613
rect 50 -75637 108 -75625
rect 50 -76613 62 -75637
rect 96 -76613 108 -75637
rect 50 -76625 108 -76613
rect -108 -76855 -50 -76843
rect -108 -77831 -96 -76855
rect -62 -77831 -50 -76855
rect -108 -77843 -50 -77831
rect 50 -76855 108 -76843
rect 50 -77831 62 -76855
rect 96 -77831 108 -76855
rect 50 -77843 108 -77831
rect -108 -78073 -50 -78061
rect -108 -79049 -96 -78073
rect -62 -79049 -50 -78073
rect -108 -79061 -50 -79049
rect 50 -78073 108 -78061
rect 50 -79049 62 -78073
rect 96 -79049 108 -78073
rect 50 -79061 108 -79049
rect -108 -79291 -50 -79279
rect -108 -80267 -96 -79291
rect -62 -80267 -50 -79291
rect -108 -80279 -50 -80267
rect 50 -79291 108 -79279
rect 50 -80267 62 -79291
rect 96 -80267 108 -79291
rect 50 -80279 108 -80267
rect -108 -80509 -50 -80497
rect -108 -81485 -96 -80509
rect -62 -81485 -50 -80509
rect -108 -81497 -50 -81485
rect 50 -80509 108 -80497
rect 50 -81485 62 -80509
rect 96 -81485 108 -80509
rect 50 -81497 108 -81485
rect -108 -81727 -50 -81715
rect -108 -82703 -96 -81727
rect -62 -82703 -50 -81727
rect -108 -82715 -50 -82703
rect 50 -81727 108 -81715
rect 50 -82703 62 -81727
rect 96 -82703 108 -81727
rect 50 -82715 108 -82703
rect -108 -82945 -50 -82933
rect -108 -83921 -96 -82945
rect -62 -83921 -50 -82945
rect -108 -83933 -50 -83921
rect 50 -82945 108 -82933
rect 50 -83921 62 -82945
rect 96 -83921 108 -82945
rect 50 -83933 108 -83921
rect -108 -84163 -50 -84151
rect -108 -85139 -96 -84163
rect -62 -85139 -50 -84163
rect -108 -85151 -50 -85139
rect 50 -84163 108 -84151
rect 50 -85139 62 -84163
rect 96 -85139 108 -84163
rect 50 -85151 108 -85139
rect -108 -85381 -50 -85369
rect -108 -86357 -96 -85381
rect -62 -86357 -50 -85381
rect -108 -86369 -50 -86357
rect 50 -85381 108 -85369
rect 50 -86357 62 -85381
rect 96 -86357 108 -85381
rect 50 -86369 108 -86357
rect -108 -86599 -50 -86587
rect -108 -87575 -96 -86599
rect -62 -87575 -50 -86599
rect -108 -87587 -50 -87575
rect 50 -86599 108 -86587
rect 50 -87575 62 -86599
rect 96 -87575 108 -86599
rect 50 -87587 108 -87575
rect -108 -87817 -50 -87805
rect -108 -88793 -96 -87817
rect -62 -88793 -50 -87817
rect -108 -88805 -50 -88793
rect 50 -87817 108 -87805
rect 50 -88793 62 -87817
rect 96 -88793 108 -87817
rect 50 -88805 108 -88793
rect -108 -89035 -50 -89023
rect -108 -90011 -96 -89035
rect -62 -90011 -50 -89035
rect -108 -90023 -50 -90011
rect 50 -89035 108 -89023
rect 50 -90011 62 -89035
rect 96 -90011 108 -89035
rect 50 -90023 108 -90011
rect -108 -90253 -50 -90241
rect -108 -91229 -96 -90253
rect -62 -91229 -50 -90253
rect -108 -91241 -50 -91229
rect 50 -90253 108 -90241
rect 50 -91229 62 -90253
rect 96 -91229 108 -90253
rect 50 -91241 108 -91229
rect -108 -91471 -50 -91459
rect -108 -92447 -96 -91471
rect -62 -92447 -50 -91471
rect -108 -92459 -50 -92447
rect 50 -91471 108 -91459
rect 50 -92447 62 -91471
rect 96 -92447 108 -91471
rect 50 -92459 108 -92447
rect -108 -92689 -50 -92677
rect -108 -93665 -96 -92689
rect -62 -93665 -50 -92689
rect -108 -93677 -50 -93665
rect 50 -92689 108 -92677
rect 50 -93665 62 -92689
rect 96 -93665 108 -92689
rect 50 -93677 108 -93665
rect -108 -93907 -50 -93895
rect -108 -94883 -96 -93907
rect -62 -94883 -50 -93907
rect -108 -94895 -50 -94883
rect 50 -93907 108 -93895
rect 50 -94883 62 -93907
rect 96 -94883 108 -93907
rect 50 -94895 108 -94883
rect -108 -95125 -50 -95113
rect -108 -96101 -96 -95125
rect -62 -96101 -50 -95125
rect -108 -96113 -50 -96101
rect 50 -95125 108 -95113
rect 50 -96101 62 -95125
rect 96 -96101 108 -95125
rect 50 -96113 108 -96101
rect -108 -96343 -50 -96331
rect -108 -97319 -96 -96343
rect -62 -97319 -50 -96343
rect -108 -97331 -50 -97319
rect 50 -96343 108 -96331
rect 50 -97319 62 -96343
rect 96 -97319 108 -96343
rect 50 -97331 108 -97319
rect -108 -97561 -50 -97549
rect -108 -98537 -96 -97561
rect -62 -98537 -50 -97561
rect -108 -98549 -50 -98537
rect 50 -97561 108 -97549
rect 50 -98537 62 -97561
rect 96 -98537 108 -97561
rect 50 -98549 108 -98537
rect -108 -98779 -50 -98767
rect -108 -99755 -96 -98779
rect -62 -99755 -50 -98779
rect -108 -99767 -50 -99755
rect 50 -98779 108 -98767
rect 50 -99755 62 -98779
rect 96 -99755 108 -98779
rect 50 -99767 108 -99755
rect -108 -99997 -50 -99985
rect -108 -100973 -96 -99997
rect -62 -100973 -50 -99997
rect -108 -100985 -50 -100973
rect 50 -99997 108 -99985
rect 50 -100973 62 -99997
rect 96 -100973 108 -99997
rect 50 -100985 108 -100973
rect -108 -101215 -50 -101203
rect -108 -102191 -96 -101215
rect -62 -102191 -50 -101215
rect -108 -102203 -50 -102191
rect 50 -101215 108 -101203
rect 50 -102191 62 -101215
rect 96 -102191 108 -101215
rect 50 -102203 108 -102191
rect -108 -102433 -50 -102421
rect -108 -103409 -96 -102433
rect -62 -103409 -50 -102433
rect -108 -103421 -50 -103409
rect 50 -102433 108 -102421
rect 50 -103409 62 -102433
rect 96 -103409 108 -102433
rect 50 -103421 108 -103409
rect -108 -103651 -50 -103639
rect -108 -104627 -96 -103651
rect -62 -104627 -50 -103651
rect -108 -104639 -50 -104627
rect 50 -103651 108 -103639
rect 50 -104627 62 -103651
rect 96 -104627 108 -103651
rect 50 -104639 108 -104627
rect -108 -104869 -50 -104857
rect -108 -105845 -96 -104869
rect -62 -105845 -50 -104869
rect -108 -105857 -50 -105845
rect 50 -104869 108 -104857
rect 50 -105845 62 -104869
rect 96 -105845 108 -104869
rect 50 -105857 108 -105845
rect -108 -106087 -50 -106075
rect -108 -107063 -96 -106087
rect -62 -107063 -50 -106087
rect -108 -107075 -50 -107063
rect 50 -106087 108 -106075
rect 50 -107063 62 -106087
rect 96 -107063 108 -106087
rect 50 -107075 108 -107063
rect -108 -107305 -50 -107293
rect -108 -108281 -96 -107305
rect -62 -108281 -50 -107305
rect -108 -108293 -50 -108281
rect 50 -107305 108 -107293
rect 50 -108281 62 -107305
rect 96 -108281 108 -107305
rect 50 -108293 108 -108281
rect -108 -108523 -50 -108511
rect -108 -109499 -96 -108523
rect -62 -109499 -50 -108523
rect -108 -109511 -50 -109499
rect 50 -108523 108 -108511
rect 50 -109499 62 -108523
rect 96 -109499 108 -108523
rect 50 -109511 108 -109499
rect -108 -109741 -50 -109729
rect -108 -110717 -96 -109741
rect -62 -110717 -50 -109741
rect -108 -110729 -50 -110717
rect 50 -109741 108 -109729
rect 50 -110717 62 -109741
rect 96 -110717 108 -109741
rect 50 -110729 108 -110717
rect -108 -110959 -50 -110947
rect -108 -111935 -96 -110959
rect -62 -111935 -50 -110959
rect -108 -111947 -50 -111935
rect 50 -110959 108 -110947
rect 50 -111935 62 -110959
rect 96 -111935 108 -110959
rect 50 -111947 108 -111935
rect -108 -112177 -50 -112165
rect -108 -113153 -96 -112177
rect -62 -113153 -50 -112177
rect -108 -113165 -50 -113153
rect 50 -112177 108 -112165
rect 50 -113153 62 -112177
rect 96 -113153 108 -112177
rect 50 -113165 108 -113153
rect -108 -113395 -50 -113383
rect -108 -114371 -96 -113395
rect -62 -114371 -50 -113395
rect -108 -114383 -50 -114371
rect 50 -113395 108 -113383
rect 50 -114371 62 -113395
rect 96 -114371 108 -113395
rect 50 -114383 108 -114371
rect -108 -114613 -50 -114601
rect -108 -115589 -96 -114613
rect -62 -115589 -50 -114613
rect -108 -115601 -50 -115589
rect 50 -114613 108 -114601
rect 50 -115589 62 -114613
rect 96 -115589 108 -114613
rect 50 -115601 108 -115589
rect -108 -115831 -50 -115819
rect -108 -116807 -96 -115831
rect -62 -116807 -50 -115831
rect -108 -116819 -50 -116807
rect 50 -115831 108 -115819
rect 50 -116807 62 -115831
rect 96 -116807 108 -115831
rect 50 -116819 108 -116807
rect -108 -117049 -50 -117037
rect -108 -118025 -96 -117049
rect -62 -118025 -50 -117049
rect -108 -118037 -50 -118025
rect 50 -117049 108 -117037
rect 50 -118025 62 -117049
rect 96 -118025 108 -117049
rect 50 -118037 108 -118025
rect -108 -118267 -50 -118255
rect -108 -119243 -96 -118267
rect -62 -119243 -50 -118267
rect -108 -119255 -50 -119243
rect 50 -118267 108 -118255
rect 50 -119243 62 -118267
rect 96 -119243 108 -118267
rect 50 -119255 108 -119243
rect -108 -119485 -50 -119473
rect -108 -120461 -96 -119485
rect -62 -120461 -50 -119485
rect -108 -120473 -50 -120461
rect 50 -119485 108 -119473
rect 50 -120461 62 -119485
rect 96 -120461 108 -119485
rect 50 -120473 108 -120461
rect -108 -120703 -50 -120691
rect -108 -121679 -96 -120703
rect -62 -121679 -50 -120703
rect -108 -121691 -50 -121679
rect 50 -120703 108 -120691
rect 50 -121679 62 -120703
rect 96 -121679 108 -120703
rect 50 -121691 108 -121679
rect -108 -121921 -50 -121909
rect -108 -122897 -96 -121921
rect -62 -122897 -50 -121921
rect -108 -122909 -50 -122897
rect 50 -121921 108 -121909
rect 50 -122897 62 -121921
rect 96 -122897 108 -121921
rect 50 -122909 108 -122897
rect -108 -123139 -50 -123127
rect -108 -124115 -96 -123139
rect -62 -124115 -50 -123139
rect -108 -124127 -50 -124115
rect 50 -123139 108 -123127
rect 50 -124115 62 -123139
rect 96 -124115 108 -123139
rect 50 -124127 108 -124115
rect -108 -124357 -50 -124345
rect -108 -125333 -96 -124357
rect -62 -125333 -50 -124357
rect -108 -125345 -50 -125333
rect 50 -124357 108 -124345
rect 50 -125333 62 -124357
rect 96 -125333 108 -124357
rect 50 -125345 108 -125333
rect -108 -125575 -50 -125563
rect -108 -126551 -96 -125575
rect -62 -126551 -50 -125575
rect -108 -126563 -50 -126551
rect 50 -125575 108 -125563
rect 50 -126551 62 -125575
rect 96 -126551 108 -125575
rect 50 -126563 108 -126551
rect -108 -126793 -50 -126781
rect -108 -127769 -96 -126793
rect -62 -127769 -50 -126793
rect -108 -127781 -50 -127769
rect 50 -126793 108 -126781
rect 50 -127769 62 -126793
rect 96 -127769 108 -126793
rect 50 -127781 108 -127769
rect -108 -128011 -50 -127999
rect -108 -128987 -96 -128011
rect -62 -128987 -50 -128011
rect -108 -128999 -50 -128987
rect 50 -128011 108 -127999
rect 50 -128987 62 -128011
rect 96 -128987 108 -128011
rect 50 -128999 108 -128987
rect -108 -129229 -50 -129217
rect -108 -130205 -96 -129229
rect -62 -130205 -50 -129229
rect -108 -130217 -50 -130205
rect 50 -129229 108 -129217
rect 50 -130205 62 -129229
rect 96 -130205 108 -129229
rect 50 -130217 108 -130205
rect -108 -130447 -50 -130435
rect -108 -131423 -96 -130447
rect -62 -131423 -50 -130447
rect -108 -131435 -50 -131423
rect 50 -130447 108 -130435
rect 50 -131423 62 -130447
rect 96 -131423 108 -130447
rect 50 -131435 108 -131423
rect -108 -131665 -50 -131653
rect -108 -132641 -96 -131665
rect -62 -132641 -50 -131665
rect -108 -132653 -50 -132641
rect 50 -131665 108 -131653
rect 50 -132641 62 -131665
rect 96 -132641 108 -131665
rect 50 -132653 108 -132641
rect -108 -132883 -50 -132871
rect -108 -133859 -96 -132883
rect -62 -133859 -50 -132883
rect -108 -133871 -50 -133859
rect 50 -132883 108 -132871
rect 50 -133859 62 -132883
rect 96 -133859 108 -132883
rect 50 -133871 108 -133859
rect -108 -134101 -50 -134089
rect -108 -135077 -96 -134101
rect -62 -135077 -50 -134101
rect -108 -135089 -50 -135077
rect 50 -134101 108 -134089
rect 50 -135077 62 -134101
rect 96 -135077 108 -134101
rect 50 -135089 108 -135077
rect -108 -135319 -50 -135307
rect -108 -136295 -96 -135319
rect -62 -136295 -50 -135319
rect -108 -136307 -50 -136295
rect 50 -135319 108 -135307
rect 50 -136295 62 -135319
rect 96 -136295 108 -135319
rect 50 -136307 108 -136295
rect -108 -136537 -50 -136525
rect -108 -137513 -96 -136537
rect -62 -137513 -50 -136537
rect -108 -137525 -50 -137513
rect 50 -136537 108 -136525
rect 50 -137513 62 -136537
rect 96 -137513 108 -136537
rect 50 -137525 108 -137513
rect -108 -137755 -50 -137743
rect -108 -138731 -96 -137755
rect -62 -138731 -50 -137755
rect -108 -138743 -50 -138731
rect 50 -137755 108 -137743
rect 50 -138731 62 -137755
rect 96 -138731 108 -137755
rect 50 -138743 108 -138731
rect -108 -138973 -50 -138961
rect -108 -139949 -96 -138973
rect -62 -139949 -50 -138973
rect -108 -139961 -50 -139949
rect 50 -138973 108 -138961
rect 50 -139949 62 -138973
rect 96 -139949 108 -138973
rect 50 -139961 108 -139949
rect -108 -140191 -50 -140179
rect -108 -141167 -96 -140191
rect -62 -141167 -50 -140191
rect -108 -141179 -50 -141167
rect 50 -140191 108 -140179
rect 50 -141167 62 -140191
rect 96 -141167 108 -140191
rect 50 -141179 108 -141167
rect -108 -141409 -50 -141397
rect -108 -142385 -96 -141409
rect -62 -142385 -50 -141409
rect -108 -142397 -50 -142385
rect 50 -141409 108 -141397
rect 50 -142385 62 -141409
rect 96 -142385 108 -141409
rect 50 -142397 108 -142385
rect -108 -142627 -50 -142615
rect -108 -143603 -96 -142627
rect -62 -143603 -50 -142627
rect -108 -143615 -50 -143603
rect 50 -142627 108 -142615
rect 50 -143603 62 -142627
rect 96 -143603 108 -142627
rect 50 -143615 108 -143603
rect -108 -143845 -50 -143833
rect -108 -144821 -96 -143845
rect -62 -144821 -50 -143845
rect -108 -144833 -50 -144821
rect 50 -143845 108 -143833
rect 50 -144821 62 -143845
rect 96 -144821 108 -143845
rect 50 -144833 108 -144821
rect -108 -145063 -50 -145051
rect -108 -146039 -96 -145063
rect -62 -146039 -50 -145063
rect -108 -146051 -50 -146039
rect 50 -145063 108 -145051
rect 50 -146039 62 -145063
rect 96 -146039 108 -145063
rect 50 -146051 108 -146039
rect -108 -146281 -50 -146269
rect -108 -147257 -96 -146281
rect -62 -147257 -50 -146281
rect -108 -147269 -50 -147257
rect 50 -146281 108 -146269
rect 50 -147257 62 -146281
rect 96 -147257 108 -146281
rect 50 -147269 108 -147257
rect -108 -147499 -50 -147487
rect -108 -148475 -96 -147499
rect -62 -148475 -50 -147499
rect -108 -148487 -50 -148475
rect 50 -147499 108 -147487
rect 50 -148475 62 -147499
rect 96 -148475 108 -147499
rect 50 -148487 108 -148475
rect -108 -148717 -50 -148705
rect -108 -149693 -96 -148717
rect -62 -149693 -50 -148717
rect -108 -149705 -50 -149693
rect 50 -148717 108 -148705
rect 50 -149693 62 -148717
rect 96 -149693 108 -148717
rect 50 -149705 108 -149693
rect -108 -149935 -50 -149923
rect -108 -150911 -96 -149935
rect -62 -150911 -50 -149935
rect -108 -150923 -50 -150911
rect 50 -149935 108 -149923
rect 50 -150911 62 -149935
rect 96 -150911 108 -149935
rect 50 -150923 108 -150911
rect -108 -151153 -50 -151141
rect -108 -152129 -96 -151153
rect -62 -152129 -50 -151153
rect -108 -152141 -50 -152129
rect 50 -151153 108 -151141
rect 50 -152129 62 -151153
rect 96 -152129 108 -151153
rect 50 -152141 108 -152129
rect -108 -152371 -50 -152359
rect -108 -153347 -96 -152371
rect -62 -153347 -50 -152371
rect -108 -153359 -50 -153347
rect 50 -152371 108 -152359
rect 50 -153347 62 -152371
rect 96 -153347 108 -152371
rect 50 -153359 108 -153347
rect -108 -153589 -50 -153577
rect -108 -154565 -96 -153589
rect -62 -154565 -50 -153589
rect -108 -154577 -50 -154565
rect 50 -153589 108 -153577
rect 50 -154565 62 -153589
rect 96 -154565 108 -153589
rect 50 -154577 108 -154565
rect -108 -154807 -50 -154795
rect -108 -155783 -96 -154807
rect -62 -155783 -50 -154807
rect -108 -155795 -50 -155783
rect 50 -154807 108 -154795
rect 50 -155783 62 -154807
rect 96 -155783 108 -154807
rect 50 -155795 108 -155783
rect -108 -156025 -50 -156013
rect -108 -157001 -96 -156025
rect -62 -157001 -50 -156025
rect -108 -157013 -50 -157001
rect 50 -156025 108 -156013
rect 50 -157001 62 -156025
rect 96 -157001 108 -156025
rect 50 -157013 108 -157001
rect -108 -157243 -50 -157231
rect -108 -158219 -96 -157243
rect -62 -158219 -50 -157243
rect -108 -158231 -50 -158219
rect 50 -157243 108 -157231
rect 50 -158219 62 -157243
rect 96 -158219 108 -157243
rect 50 -158231 108 -158219
rect -108 -158461 -50 -158449
rect -108 -159437 -96 -158461
rect -62 -159437 -50 -158461
rect -108 -159449 -50 -159437
rect 50 -158461 108 -158449
rect 50 -159437 62 -158461
rect 96 -159437 108 -158461
rect 50 -159449 108 -159437
rect -108 -159679 -50 -159667
rect -108 -160655 -96 -159679
rect -62 -160655 -50 -159679
rect -108 -160667 -50 -160655
rect 50 -159679 108 -159667
rect 50 -160655 62 -159679
rect 96 -160655 108 -159679
rect 50 -160667 108 -160655
rect -108 -160897 -50 -160885
rect -108 -161873 -96 -160897
rect -62 -161873 -50 -160897
rect -108 -161885 -50 -161873
rect 50 -160897 108 -160885
rect 50 -161873 62 -160897
rect 96 -161873 108 -160897
rect 50 -161885 108 -161873
rect -108 -162115 -50 -162103
rect -108 -163091 -96 -162115
rect -62 -163091 -50 -162115
rect -108 -163103 -50 -163091
rect 50 -162115 108 -162103
rect 50 -163091 62 -162115
rect 96 -163091 108 -162115
rect 50 -163103 108 -163091
rect -108 -163333 -50 -163321
rect -108 -164309 -96 -163333
rect -62 -164309 -50 -163333
rect -108 -164321 -50 -164309
rect 50 -163333 108 -163321
rect 50 -164309 62 -163333
rect 96 -164309 108 -163333
rect 50 -164321 108 -164309
rect -108 -164551 -50 -164539
rect -108 -165527 -96 -164551
rect -62 -165527 -50 -164551
rect -108 -165539 -50 -165527
rect 50 -164551 108 -164539
rect 50 -165527 62 -164551
rect 96 -165527 108 -164551
rect 50 -165539 108 -165527
rect -108 -165769 -50 -165757
rect -108 -166745 -96 -165769
rect -62 -166745 -50 -165769
rect -108 -166757 -50 -166745
rect 50 -165769 108 -165757
rect 50 -166745 62 -165769
rect 96 -166745 108 -165769
rect 50 -166757 108 -166745
rect -108 -166987 -50 -166975
rect -108 -167963 -96 -166987
rect -62 -167963 -50 -166987
rect -108 -167975 -50 -167963
rect 50 -166987 108 -166975
rect 50 -167963 62 -166987
rect 96 -167963 108 -166987
rect 50 -167975 108 -167963
rect -108 -168205 -50 -168193
rect -108 -169181 -96 -168205
rect -62 -169181 -50 -168205
rect -108 -169193 -50 -169181
rect 50 -168205 108 -168193
rect 50 -169181 62 -168205
rect 96 -169181 108 -168205
rect 50 -169193 108 -169181
rect -108 -169423 -50 -169411
rect -108 -170399 -96 -169423
rect -62 -170399 -50 -169423
rect -108 -170411 -50 -170399
rect 50 -169423 108 -169411
rect 50 -170399 62 -169423
rect 96 -170399 108 -169423
rect 50 -170411 108 -170399
rect -108 -170641 -50 -170629
rect -108 -171617 -96 -170641
rect -62 -171617 -50 -170641
rect -108 -171629 -50 -171617
rect 50 -170641 108 -170629
rect 50 -171617 62 -170641
rect 96 -171617 108 -170641
rect 50 -171629 108 -171617
rect -108 -171859 -50 -171847
rect -108 -172835 -96 -171859
rect -62 -172835 -50 -171859
rect -108 -172847 -50 -172835
rect 50 -171859 108 -171847
rect 50 -172835 62 -171859
rect 96 -172835 108 -171859
rect 50 -172847 108 -172835
rect -108 -173077 -50 -173065
rect -108 -174053 -96 -173077
rect -62 -174053 -50 -173077
rect -108 -174065 -50 -174053
rect 50 -173077 108 -173065
rect 50 -174053 62 -173077
rect 96 -174053 108 -173077
rect 50 -174065 108 -174053
rect -108 -174295 -50 -174283
rect -108 -175271 -96 -174295
rect -62 -175271 -50 -174295
rect -108 -175283 -50 -175271
rect 50 -174295 108 -174283
rect 50 -175271 62 -174295
rect 96 -175271 108 -174295
rect 50 -175283 108 -175271
rect -108 -175513 -50 -175501
rect -108 -176489 -96 -175513
rect -62 -176489 -50 -175513
rect -108 -176501 -50 -176489
rect 50 -175513 108 -175501
rect 50 -176489 62 -175513
rect 96 -176489 108 -175513
rect 50 -176501 108 -176489
rect -108 -176731 -50 -176719
rect -108 -177707 -96 -176731
rect -62 -177707 -50 -176731
rect -108 -177719 -50 -177707
rect 50 -176731 108 -176719
rect 50 -177707 62 -176731
rect 96 -177707 108 -176731
rect 50 -177719 108 -177707
rect -108 -177949 -50 -177937
rect -108 -178925 -96 -177949
rect -62 -178925 -50 -177949
rect -108 -178937 -50 -178925
rect 50 -177949 108 -177937
rect 50 -178925 62 -177949
rect 96 -178925 108 -177949
rect 50 -178937 108 -178925
rect -108 -179167 -50 -179155
rect -108 -180143 -96 -179167
rect -62 -180143 -50 -179167
rect -108 -180155 -50 -180143
rect 50 -179167 108 -179155
rect 50 -180143 62 -179167
rect 96 -180143 108 -179167
rect 50 -180155 108 -180143
rect -108 -180385 -50 -180373
rect -108 -181361 -96 -180385
rect -62 -181361 -50 -180385
rect -108 -181373 -50 -181361
rect 50 -180385 108 -180373
rect 50 -181361 62 -180385
rect 96 -181361 108 -180385
rect 50 -181373 108 -181361
rect -108 -181603 -50 -181591
rect -108 -182579 -96 -181603
rect -62 -182579 -50 -181603
rect -108 -182591 -50 -182579
rect 50 -181603 108 -181591
rect 50 -182579 62 -181603
rect 96 -182579 108 -181603
rect 50 -182591 108 -182579
rect -108 -182821 -50 -182809
rect -108 -183797 -96 -182821
rect -62 -183797 -50 -182821
rect -108 -183809 -50 -183797
rect 50 -182821 108 -182809
rect 50 -183797 62 -182821
rect 96 -183797 108 -182821
rect 50 -183809 108 -183797
rect -108 -184039 -50 -184027
rect -108 -185015 -96 -184039
rect -62 -185015 -50 -184039
rect -108 -185027 -50 -185015
rect 50 -184039 108 -184027
rect 50 -185015 62 -184039
rect 96 -185015 108 -184039
rect 50 -185027 108 -185015
rect -108 -185257 -50 -185245
rect -108 -186233 -96 -185257
rect -62 -186233 -50 -185257
rect -108 -186245 -50 -186233
rect 50 -185257 108 -185245
rect 50 -186233 62 -185257
rect 96 -186233 108 -185257
rect 50 -186245 108 -186233
rect -108 -186475 -50 -186463
rect -108 -187451 -96 -186475
rect -62 -187451 -50 -186475
rect -108 -187463 -50 -187451
rect 50 -186475 108 -186463
rect 50 -187451 62 -186475
rect 96 -187451 108 -186475
rect 50 -187463 108 -187451
rect -108 -187693 -50 -187681
rect -108 -188669 -96 -187693
rect -62 -188669 -50 -187693
rect -108 -188681 -50 -188669
rect 50 -187693 108 -187681
rect 50 -188669 62 -187693
rect 96 -188669 108 -187693
rect 50 -188681 108 -188669
rect -108 -188911 -50 -188899
rect -108 -189887 -96 -188911
rect -62 -189887 -50 -188911
rect -108 -189899 -50 -189887
rect 50 -188911 108 -188899
rect 50 -189887 62 -188911
rect 96 -189887 108 -188911
rect 50 -189899 108 -189887
rect -108 -190129 -50 -190117
rect -108 -191105 -96 -190129
rect -62 -191105 -50 -190129
rect -108 -191117 -50 -191105
rect 50 -190129 108 -190117
rect 50 -191105 62 -190129
rect 96 -191105 108 -190129
rect 50 -191117 108 -191105
rect -108 -191347 -50 -191335
rect -108 -192323 -96 -191347
rect -62 -192323 -50 -191347
rect -108 -192335 -50 -192323
rect 50 -191347 108 -191335
rect 50 -192323 62 -191347
rect 96 -192323 108 -191347
rect 50 -192335 108 -192323
rect -108 -192565 -50 -192553
rect -108 -193541 -96 -192565
rect -62 -193541 -50 -192565
rect -108 -193553 -50 -193541
rect 50 -192565 108 -192553
rect 50 -193541 62 -192565
rect 96 -193541 108 -192565
rect 50 -193553 108 -193541
rect -108 -193783 -50 -193771
rect -108 -194759 -96 -193783
rect -62 -194759 -50 -193783
rect -108 -194771 -50 -194759
rect 50 -193783 108 -193771
rect 50 -194759 62 -193783
rect 96 -194759 108 -193783
rect 50 -194771 108 -194759
rect -108 -195001 -50 -194989
rect -108 -195977 -96 -195001
rect -62 -195977 -50 -195001
rect -108 -195989 -50 -195977
rect 50 -195001 108 -194989
rect 50 -195977 62 -195001
rect 96 -195977 108 -195001
rect 50 -195989 108 -195977
rect -108 -196219 -50 -196207
rect -108 -197195 -96 -196219
rect -62 -197195 -50 -196219
rect -108 -197207 -50 -197195
rect 50 -196219 108 -196207
rect 50 -197195 62 -196219
rect 96 -197195 108 -196219
rect 50 -197207 108 -197195
rect -108 -197437 -50 -197425
rect -108 -198413 -96 -197437
rect -62 -198413 -50 -197437
rect -108 -198425 -50 -198413
rect 50 -197437 108 -197425
rect 50 -198413 62 -197437
rect 96 -198413 108 -197437
rect 50 -198425 108 -198413
rect -108 -198655 -50 -198643
rect -108 -199631 -96 -198655
rect -62 -199631 -50 -198655
rect -108 -199643 -50 -199631
rect 50 -198655 108 -198643
rect 50 -199631 62 -198655
rect 96 -199631 108 -198655
rect 50 -199643 108 -199631
rect -108 -199873 -50 -199861
rect -108 -200849 -96 -199873
rect -62 -200849 -50 -199873
rect -108 -200861 -50 -200849
rect 50 -199873 108 -199861
rect 50 -200849 62 -199873
rect 96 -200849 108 -199873
rect 50 -200861 108 -200849
rect -108 -201091 -50 -201079
rect -108 -202067 -96 -201091
rect -62 -202067 -50 -201091
rect -108 -202079 -50 -202067
rect 50 -201091 108 -201079
rect 50 -202067 62 -201091
rect 96 -202067 108 -201091
rect 50 -202079 108 -202067
rect -108 -202309 -50 -202297
rect -108 -203285 -96 -202309
rect -62 -203285 -50 -202309
rect -108 -203297 -50 -203285
rect 50 -202309 108 -202297
rect 50 -203285 62 -202309
rect 96 -203285 108 -202309
rect 50 -203297 108 -203285
rect -108 -203527 -50 -203515
rect -108 -204503 -96 -203527
rect -62 -204503 -50 -203527
rect -108 -204515 -50 -204503
rect 50 -203527 108 -203515
rect 50 -204503 62 -203527
rect 96 -204503 108 -203527
rect 50 -204515 108 -204503
rect -108 -204745 -50 -204733
rect -108 -205721 -96 -204745
rect -62 -205721 -50 -204745
rect -108 -205733 -50 -205721
rect 50 -204745 108 -204733
rect 50 -205721 62 -204745
rect 96 -205721 108 -204745
rect 50 -205733 108 -205721
rect -108 -205963 -50 -205951
rect -108 -206939 -96 -205963
rect -62 -206939 -50 -205963
rect -108 -206951 -50 -206939
rect 50 -205963 108 -205951
rect 50 -206939 62 -205963
rect 96 -206939 108 -205963
rect 50 -206951 108 -206939
rect -108 -207181 -50 -207169
rect -108 -208157 -96 -207181
rect -62 -208157 -50 -207181
rect -108 -208169 -50 -208157
rect 50 -207181 108 -207169
rect 50 -208157 62 -207181
rect 96 -208157 108 -207181
rect 50 -208169 108 -208157
rect -108 -208399 -50 -208387
rect -108 -209375 -96 -208399
rect -62 -209375 -50 -208399
rect -108 -209387 -50 -209375
rect 50 -208399 108 -208387
rect 50 -209375 62 -208399
rect 96 -209375 108 -208399
rect 50 -209387 108 -209375
rect -108 -209617 -50 -209605
rect -108 -210593 -96 -209617
rect -62 -210593 -50 -209617
rect -108 -210605 -50 -210593
rect 50 -209617 108 -209605
rect 50 -210593 62 -209617
rect 96 -210593 108 -209617
rect 50 -210605 108 -210593
rect -108 -210835 -50 -210823
rect -108 -211811 -96 -210835
rect -62 -211811 -50 -210835
rect -108 -211823 -50 -211811
rect 50 -210835 108 -210823
rect 50 -211811 62 -210835
rect 96 -211811 108 -210835
rect 50 -211823 108 -211811
rect -108 -212053 -50 -212041
rect -108 -213029 -96 -212053
rect -62 -213029 -50 -212053
rect -108 -213041 -50 -213029
rect 50 -212053 108 -212041
rect 50 -213029 62 -212053
rect 96 -213029 108 -212053
rect 50 -213041 108 -213029
rect -108 -213271 -50 -213259
rect -108 -214247 -96 -213271
rect -62 -214247 -50 -213271
rect -108 -214259 -50 -214247
rect 50 -213271 108 -213259
rect 50 -214247 62 -213271
rect 96 -214247 108 -213271
rect 50 -214259 108 -214247
rect -108 -214489 -50 -214477
rect -108 -215465 -96 -214489
rect -62 -215465 -50 -214489
rect -108 -215477 -50 -215465
rect 50 -214489 108 -214477
rect 50 -215465 62 -214489
rect 96 -215465 108 -214489
rect 50 -215477 108 -215465
rect -108 -215707 -50 -215695
rect -108 -216683 -96 -215707
rect -62 -216683 -50 -215707
rect -108 -216695 -50 -216683
rect 50 -215707 108 -215695
rect 50 -216683 62 -215707
rect 96 -216683 108 -215707
rect 50 -216695 108 -216683
rect -108 -216925 -50 -216913
rect -108 -217901 -96 -216925
rect -62 -217901 -50 -216925
rect -108 -217913 -50 -217901
rect 50 -216925 108 -216913
rect 50 -217901 62 -216925
rect 96 -217901 108 -216925
rect 50 -217913 108 -217901
rect -108 -218143 -50 -218131
rect -108 -219119 -96 -218143
rect -62 -219119 -50 -218143
rect -108 -219131 -50 -219119
rect 50 -218143 108 -218131
rect 50 -219119 62 -218143
rect 96 -219119 108 -218143
rect 50 -219131 108 -219119
rect -108 -219361 -50 -219349
rect -108 -220337 -96 -219361
rect -62 -220337 -50 -219361
rect -108 -220349 -50 -220337
rect 50 -219361 108 -219349
rect 50 -220337 62 -219361
rect 96 -220337 108 -219361
rect 50 -220349 108 -220337
rect -108 -220579 -50 -220567
rect -108 -221555 -96 -220579
rect -62 -221555 -50 -220579
rect -108 -221567 -50 -221555
rect 50 -220579 108 -220567
rect 50 -221555 62 -220579
rect 96 -221555 108 -220579
rect 50 -221567 108 -221555
rect -108 -221797 -50 -221785
rect -108 -222773 -96 -221797
rect -62 -222773 -50 -221797
rect -108 -222785 -50 -222773
rect 50 -221797 108 -221785
rect 50 -222773 62 -221797
rect 96 -222773 108 -221797
rect 50 -222785 108 -222773
rect -108 -223015 -50 -223003
rect -108 -223991 -96 -223015
rect -62 -223991 -50 -223015
rect -108 -224003 -50 -223991
rect 50 -223015 108 -223003
rect 50 -223991 62 -223015
rect 96 -223991 108 -223015
rect 50 -224003 108 -223991
rect -108 -224233 -50 -224221
rect -108 -225209 -96 -224233
rect -62 -225209 -50 -224233
rect -108 -225221 -50 -225209
rect 50 -224233 108 -224221
rect 50 -225209 62 -224233
rect 96 -225209 108 -224233
rect 50 -225221 108 -225209
rect -108 -225451 -50 -225439
rect -108 -226427 -96 -225451
rect -62 -226427 -50 -225451
rect -108 -226439 -50 -226427
rect 50 -225451 108 -225439
rect 50 -226427 62 -225451
rect 96 -226427 108 -225451
rect 50 -226439 108 -226427
rect -108 -226669 -50 -226657
rect -108 -227645 -96 -226669
rect -62 -227645 -50 -226669
rect -108 -227657 -50 -227645
rect 50 -226669 108 -226657
rect 50 -227645 62 -226669
rect 96 -227645 108 -226669
rect 50 -227657 108 -227645
rect -108 -227887 -50 -227875
rect -108 -228863 -96 -227887
rect -62 -228863 -50 -227887
rect -108 -228875 -50 -228863
rect 50 -227887 108 -227875
rect 50 -228863 62 -227887
rect 96 -228863 108 -227887
rect 50 -228875 108 -228863
rect -108 -229105 -50 -229093
rect -108 -230081 -96 -229105
rect -62 -230081 -50 -229105
rect -108 -230093 -50 -230081
rect 50 -229105 108 -229093
rect 50 -230081 62 -229105
rect 96 -230081 108 -229105
rect 50 -230093 108 -230081
rect -108 -230323 -50 -230311
rect -108 -231299 -96 -230323
rect -62 -231299 -50 -230323
rect -108 -231311 -50 -231299
rect 50 -230323 108 -230311
rect 50 -231299 62 -230323
rect 96 -231299 108 -230323
rect 50 -231311 108 -231299
rect -108 -231541 -50 -231529
rect -108 -232517 -96 -231541
rect -62 -232517 -50 -231541
rect -108 -232529 -50 -232517
rect 50 -231541 108 -231529
rect 50 -232517 62 -231541
rect 96 -232517 108 -231541
rect 50 -232529 108 -232517
rect -108 -232759 -50 -232747
rect -108 -233735 -96 -232759
rect -62 -233735 -50 -232759
rect -108 -233747 -50 -233735
rect 50 -232759 108 -232747
rect 50 -233735 62 -232759
rect 96 -233735 108 -232759
rect 50 -233747 108 -233735
rect -108 -233977 -50 -233965
rect -108 -234953 -96 -233977
rect -62 -234953 -50 -233977
rect -108 -234965 -50 -234953
rect 50 -233977 108 -233965
rect 50 -234953 62 -233977
rect 96 -234953 108 -233977
rect 50 -234965 108 -234953
rect -108 -235195 -50 -235183
rect -108 -236171 -96 -235195
rect -62 -236171 -50 -235195
rect -108 -236183 -50 -236171
rect 50 -235195 108 -235183
rect 50 -236171 62 -235195
rect 96 -236171 108 -235195
rect 50 -236183 108 -236171
rect -108 -236413 -50 -236401
rect -108 -237389 -96 -236413
rect -62 -237389 -50 -236413
rect -108 -237401 -50 -237389
rect 50 -236413 108 -236401
rect 50 -237389 62 -236413
rect 96 -237389 108 -236413
rect 50 -237401 108 -237389
rect -108 -237631 -50 -237619
rect -108 -238607 -96 -237631
rect -62 -238607 -50 -237631
rect -108 -238619 -50 -238607
rect 50 -237631 108 -237619
rect 50 -238607 62 -237631
rect 96 -238607 108 -237631
rect 50 -238619 108 -238607
rect -108 -238849 -50 -238837
rect -108 -239825 -96 -238849
rect -62 -239825 -50 -238849
rect -108 -239837 -50 -239825
rect 50 -238849 108 -238837
rect 50 -239825 62 -238849
rect 96 -239825 108 -238849
rect 50 -239837 108 -239825
rect -108 -240067 -50 -240055
rect -108 -241043 -96 -240067
rect -62 -241043 -50 -240067
rect -108 -241055 -50 -241043
rect 50 -240067 108 -240055
rect 50 -241043 62 -240067
rect 96 -241043 108 -240067
rect 50 -241055 108 -241043
rect -108 -241285 -50 -241273
rect -108 -242261 -96 -241285
rect -62 -242261 -50 -241285
rect -108 -242273 -50 -242261
rect 50 -241285 108 -241273
rect 50 -242261 62 -241285
rect 96 -242261 108 -241285
rect 50 -242273 108 -242261
rect -108 -242503 -50 -242491
rect -108 -243479 -96 -242503
rect -62 -243479 -50 -242503
rect -108 -243491 -50 -243479
rect 50 -242503 108 -242491
rect 50 -243479 62 -242503
rect 96 -243479 108 -242503
rect 50 -243491 108 -243479
rect -108 -243721 -50 -243709
rect -108 -244697 -96 -243721
rect -62 -244697 -50 -243721
rect -108 -244709 -50 -244697
rect 50 -243721 108 -243709
rect 50 -244697 62 -243721
rect 96 -244697 108 -243721
rect 50 -244709 108 -244697
rect -108 -244939 -50 -244927
rect -108 -245915 -96 -244939
rect -62 -245915 -50 -244939
rect -108 -245927 -50 -245915
rect 50 -244939 108 -244927
rect 50 -245915 62 -244939
rect 96 -245915 108 -244939
rect 50 -245927 108 -245915
rect -108 -246157 -50 -246145
rect -108 -247133 -96 -246157
rect -62 -247133 -50 -246157
rect -108 -247145 -50 -247133
rect 50 -246157 108 -246145
rect 50 -247133 62 -246157
rect 96 -247133 108 -246157
rect 50 -247145 108 -247133
rect -108 -247375 -50 -247363
rect -108 -248351 -96 -247375
rect -62 -248351 -50 -247375
rect -108 -248363 -50 -248351
rect 50 -247375 108 -247363
rect 50 -248351 62 -247375
rect 96 -248351 108 -247375
rect 50 -248363 108 -248351
rect -108 -248593 -50 -248581
rect -108 -249569 -96 -248593
rect -62 -249569 -50 -248593
rect -108 -249581 -50 -249569
rect 50 -248593 108 -248581
rect 50 -249569 62 -248593
rect 96 -249569 108 -248593
rect 50 -249581 108 -249569
rect -108 -249811 -50 -249799
rect -108 -250787 -96 -249811
rect -62 -250787 -50 -249811
rect -108 -250799 -50 -250787
rect 50 -249811 108 -249799
rect 50 -250787 62 -249811
rect 96 -250787 108 -249811
rect 50 -250799 108 -250787
rect -108 -251029 -50 -251017
rect -108 -252005 -96 -251029
rect -62 -252005 -50 -251029
rect -108 -252017 -50 -252005
rect 50 -251029 108 -251017
rect 50 -252005 62 -251029
rect 96 -252005 108 -251029
rect 50 -252017 108 -252005
rect -108 -252247 -50 -252235
rect -108 -253223 -96 -252247
rect -62 -253223 -50 -252247
rect -108 -253235 -50 -253223
rect 50 -252247 108 -252235
rect 50 -253223 62 -252247
rect 96 -253223 108 -252247
rect 50 -253235 108 -253223
rect -108 -253465 -50 -253453
rect -108 -254441 -96 -253465
rect -62 -254441 -50 -253465
rect -108 -254453 -50 -254441
rect 50 -253465 108 -253453
rect 50 -254441 62 -253465
rect 96 -254441 108 -253465
rect 50 -254453 108 -254441
rect -108 -254683 -50 -254671
rect -108 -255659 -96 -254683
rect -62 -255659 -50 -254683
rect -108 -255671 -50 -255659
rect 50 -254683 108 -254671
rect 50 -255659 62 -254683
rect 96 -255659 108 -254683
rect 50 -255671 108 -255659
rect -108 -255901 -50 -255889
rect -108 -256877 -96 -255901
rect -62 -256877 -50 -255901
rect -108 -256889 -50 -256877
rect 50 -255901 108 -255889
rect 50 -256877 62 -255901
rect 96 -256877 108 -255901
rect 50 -256889 108 -256877
rect -108 -257119 -50 -257107
rect -108 -258095 -96 -257119
rect -62 -258095 -50 -257119
rect -108 -258107 -50 -258095
rect 50 -257119 108 -257107
rect 50 -258095 62 -257119
rect 96 -258095 108 -257119
rect 50 -258107 108 -258095
rect -108 -258337 -50 -258325
rect -108 -259313 -96 -258337
rect -62 -259313 -50 -258337
rect -108 -259325 -50 -259313
rect 50 -258337 108 -258325
rect 50 -259313 62 -258337
rect 96 -259313 108 -258337
rect 50 -259325 108 -259313
rect -108 -259555 -50 -259543
rect -108 -260531 -96 -259555
rect -62 -260531 -50 -259555
rect -108 -260543 -50 -260531
rect 50 -259555 108 -259543
rect 50 -260531 62 -259555
rect 96 -260531 108 -259555
rect 50 -260543 108 -260531
rect -108 -260773 -50 -260761
rect -108 -261749 -96 -260773
rect -62 -261749 -50 -260773
rect -108 -261761 -50 -261749
rect 50 -260773 108 -260761
rect 50 -261749 62 -260773
rect 96 -261749 108 -260773
rect 50 -261761 108 -261749
rect -108 -261991 -50 -261979
rect -108 -262967 -96 -261991
rect -62 -262967 -50 -261991
rect -108 -262979 -50 -262967
rect 50 -261991 108 -261979
rect 50 -262967 62 -261991
rect 96 -262967 108 -261991
rect 50 -262979 108 -262967
rect -108 -263209 -50 -263197
rect -108 -264185 -96 -263209
rect -62 -264185 -50 -263209
rect -108 -264197 -50 -264185
rect 50 -263209 108 -263197
rect 50 -264185 62 -263209
rect 96 -264185 108 -263209
rect 50 -264197 108 -264185
rect -108 -264427 -50 -264415
rect -108 -265403 -96 -264427
rect -62 -265403 -50 -264427
rect -108 -265415 -50 -265403
rect 50 -264427 108 -264415
rect 50 -265403 62 -264427
rect 96 -265403 108 -264427
rect 50 -265415 108 -265403
rect -108 -265645 -50 -265633
rect -108 -266621 -96 -265645
rect -62 -266621 -50 -265645
rect -108 -266633 -50 -266621
rect 50 -265645 108 -265633
rect 50 -266621 62 -265645
rect 96 -266621 108 -265645
rect 50 -266633 108 -266621
rect -108 -266863 -50 -266851
rect -108 -267839 -96 -266863
rect -62 -267839 -50 -266863
rect -108 -267851 -50 -267839
rect 50 -266863 108 -266851
rect 50 -267839 62 -266863
rect 96 -267839 108 -266863
rect 50 -267851 108 -267839
rect -108 -268081 -50 -268069
rect -108 -269057 -96 -268081
rect -62 -269057 -50 -268081
rect -108 -269069 -50 -269057
rect 50 -268081 108 -268069
rect 50 -269057 62 -268081
rect 96 -269057 108 -268081
rect 50 -269069 108 -269057
rect -108 -269299 -50 -269287
rect -108 -270275 -96 -269299
rect -62 -270275 -50 -269299
rect -108 -270287 -50 -270275
rect 50 -269299 108 -269287
rect 50 -270275 62 -269299
rect 96 -270275 108 -269299
rect 50 -270287 108 -270275
rect -108 -270517 -50 -270505
rect -108 -271493 -96 -270517
rect -62 -271493 -50 -270517
rect -108 -271505 -50 -271493
rect 50 -270517 108 -270505
rect 50 -271493 62 -270517
rect 96 -271493 108 -270517
rect 50 -271505 108 -271493
rect -108 -271735 -50 -271723
rect -108 -272711 -96 -271735
rect -62 -272711 -50 -271735
rect -108 -272723 -50 -272711
rect 50 -271735 108 -271723
rect 50 -272711 62 -271735
rect 96 -272711 108 -271735
rect 50 -272723 108 -272711
rect -108 -272953 -50 -272941
rect -108 -273929 -96 -272953
rect -62 -273929 -50 -272953
rect -108 -273941 -50 -273929
rect 50 -272953 108 -272941
rect 50 -273929 62 -272953
rect 96 -273929 108 -272953
rect 50 -273941 108 -273929
rect -108 -274171 -50 -274159
rect -108 -275147 -96 -274171
rect -62 -275147 -50 -274171
rect -108 -275159 -50 -275147
rect 50 -274171 108 -274159
rect 50 -275147 62 -274171
rect 96 -275147 108 -274171
rect 50 -275159 108 -275147
rect -108 -275389 -50 -275377
rect -108 -276365 -96 -275389
rect -62 -276365 -50 -275389
rect -108 -276377 -50 -276365
rect 50 -275389 108 -275377
rect 50 -276365 62 -275389
rect 96 -276365 108 -275389
rect 50 -276377 108 -276365
rect -108 -276607 -50 -276595
rect -108 -277583 -96 -276607
rect -62 -277583 -50 -276607
rect -108 -277595 -50 -277583
rect 50 -276607 108 -276595
rect 50 -277583 62 -276607
rect 96 -277583 108 -276607
rect 50 -277595 108 -277583
rect -108 -277825 -50 -277813
rect -108 -278801 -96 -277825
rect -62 -278801 -50 -277825
rect -108 -278813 -50 -278801
rect 50 -277825 108 -277813
rect 50 -278801 62 -277825
rect 96 -278801 108 -277825
rect 50 -278813 108 -278801
rect -108 -279043 -50 -279031
rect -108 -280019 -96 -279043
rect -62 -280019 -50 -279043
rect -108 -280031 -50 -280019
rect 50 -279043 108 -279031
rect 50 -280019 62 -279043
rect 96 -280019 108 -279043
rect 50 -280031 108 -280019
rect -108 -280261 -50 -280249
rect -108 -281237 -96 -280261
rect -62 -281237 -50 -280261
rect -108 -281249 -50 -281237
rect 50 -280261 108 -280249
rect 50 -281237 62 -280261
rect 96 -281237 108 -280261
rect 50 -281249 108 -281237
rect -108 -281479 -50 -281467
rect -108 -282455 -96 -281479
rect -62 -282455 -50 -281479
rect -108 -282467 -50 -282455
rect 50 -281479 108 -281467
rect 50 -282455 62 -281479
rect 96 -282455 108 -281479
rect 50 -282467 108 -282455
rect -108 -282697 -50 -282685
rect -108 -283673 -96 -282697
rect -62 -283673 -50 -282697
rect -108 -283685 -50 -283673
rect 50 -282697 108 -282685
rect 50 -283673 62 -282697
rect 96 -283673 108 -282697
rect 50 -283685 108 -283673
rect -108 -283915 -50 -283903
rect -108 -284891 -96 -283915
rect -62 -284891 -50 -283915
rect -108 -284903 -50 -284891
rect 50 -283915 108 -283903
rect 50 -284891 62 -283915
rect 96 -284891 108 -283915
rect 50 -284903 108 -284891
rect -108 -285133 -50 -285121
rect -108 -286109 -96 -285133
rect -62 -286109 -50 -285133
rect -108 -286121 -50 -286109
rect 50 -285133 108 -285121
rect 50 -286109 62 -285133
rect 96 -286109 108 -285133
rect 50 -286121 108 -286109
rect -108 -286351 -50 -286339
rect -108 -287327 -96 -286351
rect -62 -287327 -50 -286351
rect -108 -287339 -50 -287327
rect 50 -286351 108 -286339
rect 50 -287327 62 -286351
rect 96 -287327 108 -286351
rect 50 -287339 108 -287327
rect -108 -287569 -50 -287557
rect -108 -288545 -96 -287569
rect -62 -288545 -50 -287569
rect -108 -288557 -50 -288545
rect 50 -287569 108 -287557
rect 50 -288545 62 -287569
rect 96 -288545 108 -287569
rect 50 -288557 108 -288545
rect -108 -288787 -50 -288775
rect -108 -289763 -96 -288787
rect -62 -289763 -50 -288787
rect -108 -289775 -50 -289763
rect 50 -288787 108 -288775
rect 50 -289763 62 -288787
rect 96 -289763 108 -288787
rect 50 -289775 108 -289763
rect -108 -290005 -50 -289993
rect -108 -290981 -96 -290005
rect -62 -290981 -50 -290005
rect -108 -290993 -50 -290981
rect 50 -290005 108 -289993
rect 50 -290981 62 -290005
rect 96 -290981 108 -290005
rect 50 -290993 108 -290981
rect -108 -291223 -50 -291211
rect -108 -292199 -96 -291223
rect -62 -292199 -50 -291223
rect -108 -292211 -50 -292199
rect 50 -291223 108 -291211
rect 50 -292199 62 -291223
rect 96 -292199 108 -291223
rect 50 -292211 108 -292199
rect -108 -292441 -50 -292429
rect -108 -293417 -96 -292441
rect -62 -293417 -50 -292441
rect -108 -293429 -50 -293417
rect 50 -292441 108 -292429
rect 50 -293417 62 -292441
rect 96 -293417 108 -292441
rect 50 -293429 108 -293417
rect -108 -293659 -50 -293647
rect -108 -294635 -96 -293659
rect -62 -294635 -50 -293659
rect -108 -294647 -50 -294635
rect 50 -293659 108 -293647
rect 50 -294635 62 -293659
rect 96 -294635 108 -293659
rect 50 -294647 108 -294635
rect -108 -294877 -50 -294865
rect -108 -295853 -96 -294877
rect -62 -295853 -50 -294877
rect -108 -295865 -50 -295853
rect 50 -294877 108 -294865
rect 50 -295853 62 -294877
rect 96 -295853 108 -294877
rect 50 -295865 108 -295853
rect -108 -296095 -50 -296083
rect -108 -297071 -96 -296095
rect -62 -297071 -50 -296095
rect -108 -297083 -50 -297071
rect 50 -296095 108 -296083
rect 50 -297071 62 -296095
rect 96 -297071 108 -296095
rect 50 -297083 108 -297071
rect -108 -297313 -50 -297301
rect -108 -298289 -96 -297313
rect -62 -298289 -50 -297313
rect -108 -298301 -50 -298289
rect 50 -297313 108 -297301
rect 50 -298289 62 -297313
rect 96 -298289 108 -297313
rect 50 -298301 108 -298289
rect -108 -298531 -50 -298519
rect -108 -299507 -96 -298531
rect -62 -299507 -50 -298531
rect -108 -299519 -50 -299507
rect 50 -298531 108 -298519
rect 50 -299507 62 -298531
rect 96 -299507 108 -298531
rect 50 -299519 108 -299507
rect -108 -299749 -50 -299737
rect -108 -300725 -96 -299749
rect -62 -300725 -50 -299749
rect -108 -300737 -50 -300725
rect 50 -299749 108 -299737
rect 50 -300725 62 -299749
rect 96 -300725 108 -299749
rect 50 -300737 108 -300725
rect -108 -300967 -50 -300955
rect -108 -301943 -96 -300967
rect -62 -301943 -50 -300967
rect -108 -301955 -50 -301943
rect 50 -300967 108 -300955
rect 50 -301943 62 -300967
rect 96 -301943 108 -300967
rect 50 -301955 108 -301943
rect -108 -302185 -50 -302173
rect -108 -303161 -96 -302185
rect -62 -303161 -50 -302185
rect -108 -303173 -50 -303161
rect 50 -302185 108 -302173
rect 50 -303161 62 -302185
rect 96 -303161 108 -302185
rect 50 -303173 108 -303161
rect -108 -303403 -50 -303391
rect -108 -304379 -96 -303403
rect -62 -304379 -50 -303403
rect -108 -304391 -50 -304379
rect 50 -303403 108 -303391
rect 50 -304379 62 -303403
rect 96 -304379 108 -303403
rect 50 -304391 108 -304379
rect -108 -304621 -50 -304609
rect -108 -305597 -96 -304621
rect -62 -305597 -50 -304621
rect -108 -305609 -50 -305597
rect 50 -304621 108 -304609
rect 50 -305597 62 -304621
rect 96 -305597 108 -304621
rect 50 -305609 108 -305597
rect -108 -305839 -50 -305827
rect -108 -306815 -96 -305839
rect -62 -306815 -50 -305839
rect -108 -306827 -50 -306815
rect 50 -305839 108 -305827
rect 50 -306815 62 -305839
rect 96 -306815 108 -305839
rect 50 -306827 108 -306815
rect -108 -307057 -50 -307045
rect -108 -308033 -96 -307057
rect -62 -308033 -50 -307057
rect -108 -308045 -50 -308033
rect 50 -307057 108 -307045
rect 50 -308033 62 -307057
rect 96 -308033 108 -307057
rect 50 -308045 108 -308033
rect -108 -308275 -50 -308263
rect -108 -309251 -96 -308275
rect -62 -309251 -50 -308275
rect -108 -309263 -50 -309251
rect 50 -308275 108 -308263
rect 50 -309251 62 -308275
rect 96 -309251 108 -308275
rect 50 -309263 108 -309251
rect -108 -309493 -50 -309481
rect -108 -310469 -96 -309493
rect -62 -310469 -50 -309493
rect -108 -310481 -50 -310469
rect 50 -309493 108 -309481
rect 50 -310469 62 -309493
rect 96 -310469 108 -309493
rect 50 -310481 108 -310469
rect -108 -310711 -50 -310699
rect -108 -311687 -96 -310711
rect -62 -311687 -50 -310711
rect -108 -311699 -50 -311687
rect 50 -310711 108 -310699
rect 50 -311687 62 -310711
rect 96 -311687 108 -310711
rect 50 -311699 108 -311687
rect -108 -311929 -50 -311917
rect -108 -312905 -96 -311929
rect -62 -312905 -50 -311929
rect -108 -312917 -50 -312905
rect 50 -311929 108 -311917
rect 50 -312905 62 -311929
rect 96 -312905 108 -311929
rect 50 -312917 108 -312905
rect -108 -313147 -50 -313135
rect -108 -314123 -96 -313147
rect -62 -314123 -50 -313147
rect -108 -314135 -50 -314123
rect 50 -313147 108 -313135
rect 50 -314123 62 -313147
rect 96 -314123 108 -313147
rect 50 -314135 108 -314123
rect -108 -314365 -50 -314353
rect -108 -315341 -96 -314365
rect -62 -315341 -50 -314365
rect -108 -315353 -50 -315341
rect 50 -314365 108 -314353
rect 50 -315341 62 -314365
rect 96 -315341 108 -314365
rect 50 -315353 108 -315341
rect -108 -315583 -50 -315571
rect -108 -316559 -96 -315583
rect -62 -316559 -50 -315583
rect -108 -316571 -50 -316559
rect 50 -315583 108 -315571
rect 50 -316559 62 -315583
rect 96 -316559 108 -315583
rect 50 -316571 108 -316559
rect -108 -316801 -50 -316789
rect -108 -317777 -96 -316801
rect -62 -317777 -50 -316801
rect -108 -317789 -50 -317777
rect 50 -316801 108 -316789
rect 50 -317777 62 -316801
rect 96 -317777 108 -316801
rect 50 -317789 108 -317777
rect -108 -318019 -50 -318007
rect -108 -318995 -96 -318019
rect -62 -318995 -50 -318019
rect -108 -319007 -50 -318995
rect 50 -318019 108 -318007
rect 50 -318995 62 -318019
rect 96 -318995 108 -318019
rect 50 -319007 108 -318995
rect -108 -319237 -50 -319225
rect -108 -320213 -96 -319237
rect -62 -320213 -50 -319237
rect -108 -320225 -50 -320213
rect 50 -319237 108 -319225
rect 50 -320213 62 -319237
rect 96 -320213 108 -319237
rect 50 -320225 108 -320213
rect -108 -320455 -50 -320443
rect -108 -321431 -96 -320455
rect -62 -321431 -50 -320455
rect -108 -321443 -50 -321431
rect 50 -320455 108 -320443
rect 50 -321431 62 -320455
rect 96 -321431 108 -320455
rect 50 -321443 108 -321431
rect -108 -321673 -50 -321661
rect -108 -322649 -96 -321673
rect -62 -322649 -50 -321673
rect -108 -322661 -50 -322649
rect 50 -321673 108 -321661
rect 50 -322649 62 -321673
rect 96 -322649 108 -321673
rect 50 -322661 108 -322649
rect -108 -322891 -50 -322879
rect -108 -323867 -96 -322891
rect -62 -323867 -50 -322891
rect -108 -323879 -50 -323867
rect 50 -322891 108 -322879
rect 50 -323867 62 -322891
rect 96 -323867 108 -322891
rect 50 -323879 108 -323867
rect -108 -324109 -50 -324097
rect -108 -325085 -96 -324109
rect -62 -325085 -50 -324109
rect -108 -325097 -50 -325085
rect 50 -324109 108 -324097
rect 50 -325085 62 -324109
rect 96 -325085 108 -324109
rect 50 -325097 108 -325085
rect -108 -325327 -50 -325315
rect -108 -326303 -96 -325327
rect -62 -326303 -50 -325327
rect -108 -326315 -50 -326303
rect 50 -325327 108 -325315
rect 50 -326303 62 -325327
rect 96 -326303 108 -325327
rect 50 -326315 108 -326303
rect -108 -326545 -50 -326533
rect -108 -327521 -96 -326545
rect -62 -327521 -50 -326545
rect -108 -327533 -50 -327521
rect 50 -326545 108 -326533
rect 50 -327521 62 -326545
rect 96 -327521 108 -326545
rect 50 -327533 108 -327521
rect -108 -327763 -50 -327751
rect -108 -328739 -96 -327763
rect -62 -328739 -50 -327763
rect -108 -328751 -50 -328739
rect 50 -327763 108 -327751
rect 50 -328739 62 -327763
rect 96 -328739 108 -327763
rect 50 -328751 108 -328739
rect -108 -328981 -50 -328969
rect -108 -329957 -96 -328981
rect -62 -329957 -50 -328981
rect -108 -329969 -50 -329957
rect 50 -328981 108 -328969
rect 50 -329957 62 -328981
rect 96 -329957 108 -328981
rect 50 -329969 108 -329957
rect -108 -330199 -50 -330187
rect -108 -331175 -96 -330199
rect -62 -331175 -50 -330199
rect -108 -331187 -50 -331175
rect 50 -330199 108 -330187
rect 50 -331175 62 -330199
rect 96 -331175 108 -330199
rect 50 -331187 108 -331175
rect -108 -331417 -50 -331405
rect -108 -332393 -96 -331417
rect -62 -332393 -50 -331417
rect -108 -332405 -50 -332393
rect 50 -331417 108 -331405
rect 50 -332393 62 -331417
rect 96 -332393 108 -331417
rect 50 -332405 108 -332393
rect -108 -332635 -50 -332623
rect -108 -333611 -96 -332635
rect -62 -333611 -50 -332635
rect -108 -333623 -50 -333611
rect 50 -332635 108 -332623
rect 50 -333611 62 -332635
rect 96 -333611 108 -332635
rect 50 -333623 108 -333611
rect -108 -333853 -50 -333841
rect -108 -334829 -96 -333853
rect -62 -334829 -50 -333853
rect -108 -334841 -50 -334829
rect 50 -333853 108 -333841
rect 50 -334829 62 -333853
rect 96 -334829 108 -333853
rect 50 -334841 108 -334829
rect -108 -335071 -50 -335059
rect -108 -336047 -96 -335071
rect -62 -336047 -50 -335071
rect -108 -336059 -50 -336047
rect 50 -335071 108 -335059
rect 50 -336047 62 -335071
rect 96 -336047 108 -335071
rect 50 -336059 108 -336047
rect -108 -336289 -50 -336277
rect -108 -337265 -96 -336289
rect -62 -337265 -50 -336289
rect -108 -337277 -50 -337265
rect 50 -336289 108 -336277
rect 50 -337265 62 -336289
rect 96 -337265 108 -336289
rect 50 -337277 108 -337265
rect -108 -337507 -50 -337495
rect -108 -338483 -96 -337507
rect -62 -338483 -50 -337507
rect -108 -338495 -50 -338483
rect 50 -337507 108 -337495
rect 50 -338483 62 -337507
rect 96 -338483 108 -337507
rect 50 -338495 108 -338483
rect -108 -338725 -50 -338713
rect -108 -339701 -96 -338725
rect -62 -339701 -50 -338725
rect -108 -339713 -50 -339701
rect 50 -338725 108 -338713
rect 50 -339701 62 -338725
rect 96 -339701 108 -338725
rect 50 -339713 108 -339701
rect -108 -339943 -50 -339931
rect -108 -340919 -96 -339943
rect -62 -340919 -50 -339943
rect -108 -340931 -50 -340919
rect 50 -339943 108 -339931
rect 50 -340919 62 -339943
rect 96 -340919 108 -339943
rect 50 -340931 108 -340919
rect -108 -341161 -50 -341149
rect -108 -342137 -96 -341161
rect -62 -342137 -50 -341161
rect -108 -342149 -50 -342137
rect 50 -341161 108 -341149
rect 50 -342137 62 -341161
rect 96 -342137 108 -341161
rect 50 -342149 108 -342137
rect -108 -342379 -50 -342367
rect -108 -343355 -96 -342379
rect -62 -343355 -50 -342379
rect -108 -343367 -50 -343355
rect 50 -342379 108 -342367
rect 50 -343355 62 -342379
rect 96 -343355 108 -342379
rect 50 -343367 108 -343355
rect -108 -343597 -50 -343585
rect -108 -344573 -96 -343597
rect -62 -344573 -50 -343597
rect -108 -344585 -50 -344573
rect 50 -343597 108 -343585
rect 50 -344573 62 -343597
rect 96 -344573 108 -343597
rect 50 -344585 108 -344573
rect -108 -344815 -50 -344803
rect -108 -345791 -96 -344815
rect -62 -345791 -50 -344815
rect -108 -345803 -50 -345791
rect 50 -344815 108 -344803
rect 50 -345791 62 -344815
rect 96 -345791 108 -344815
rect 50 -345803 108 -345791
rect -108 -346033 -50 -346021
rect -108 -347009 -96 -346033
rect -62 -347009 -50 -346033
rect -108 -347021 -50 -347009
rect 50 -346033 108 -346021
rect 50 -347009 62 -346033
rect 96 -347009 108 -346033
rect 50 -347021 108 -347009
rect -108 -347251 -50 -347239
rect -108 -348227 -96 -347251
rect -62 -348227 -50 -347251
rect -108 -348239 -50 -348227
rect 50 -347251 108 -347239
rect 50 -348227 62 -347251
rect 96 -348227 108 -347251
rect 50 -348239 108 -348227
rect -108 -348469 -50 -348457
rect -108 -349445 -96 -348469
rect -62 -349445 -50 -348469
rect -108 -349457 -50 -349445
rect 50 -348469 108 -348457
rect 50 -349445 62 -348469
rect 96 -349445 108 -348469
rect 50 -349457 108 -349445
rect -108 -349687 -50 -349675
rect -108 -350663 -96 -349687
rect -62 -350663 -50 -349687
rect -108 -350675 -50 -350663
rect 50 -349687 108 -349675
rect 50 -350663 62 -349687
rect 96 -350663 108 -349687
rect 50 -350675 108 -350663
rect -108 -350905 -50 -350893
rect -108 -351881 -96 -350905
rect -62 -351881 -50 -350905
rect -108 -351893 -50 -351881
rect 50 -350905 108 -350893
rect 50 -351881 62 -350905
rect 96 -351881 108 -350905
rect 50 -351893 108 -351881
rect -108 -352123 -50 -352111
rect -108 -353099 -96 -352123
rect -62 -353099 -50 -352123
rect -108 -353111 -50 -353099
rect 50 -352123 108 -352111
rect 50 -353099 62 -352123
rect 96 -353099 108 -352123
rect 50 -353111 108 -353099
rect -108 -353341 -50 -353329
rect -108 -354317 -96 -353341
rect -62 -354317 -50 -353341
rect -108 -354329 -50 -354317
rect 50 -353341 108 -353329
rect 50 -354317 62 -353341
rect 96 -354317 108 -353341
rect 50 -354329 108 -354317
rect -108 -354559 -50 -354547
rect -108 -355535 -96 -354559
rect -62 -355535 -50 -354559
rect -108 -355547 -50 -355535
rect 50 -354559 108 -354547
rect 50 -355535 62 -354559
rect 96 -355535 108 -354559
rect 50 -355547 108 -355535
rect -108 -355777 -50 -355765
rect -108 -356753 -96 -355777
rect -62 -356753 -50 -355777
rect -108 -356765 -50 -356753
rect 50 -355777 108 -355765
rect 50 -356753 62 -355777
rect 96 -356753 108 -355777
rect 50 -356765 108 -356753
rect -108 -356995 -50 -356983
rect -108 -357971 -96 -356995
rect -62 -357971 -50 -356995
rect -108 -357983 -50 -357971
rect 50 -356995 108 -356983
rect 50 -357971 62 -356995
rect 96 -357971 108 -356995
rect 50 -357983 108 -357971
rect -108 -358213 -50 -358201
rect -108 -359189 -96 -358213
rect -62 -359189 -50 -358213
rect -108 -359201 -50 -359189
rect 50 -358213 108 -358201
rect 50 -359189 62 -358213
rect 96 -359189 108 -358213
rect 50 -359201 108 -359189
rect -108 -359431 -50 -359419
rect -108 -360407 -96 -359431
rect -62 -360407 -50 -359431
rect -108 -360419 -50 -360407
rect 50 -359431 108 -359419
rect 50 -360407 62 -359431
rect 96 -360407 108 -359431
rect 50 -360419 108 -360407
rect -108 -360649 -50 -360637
rect -108 -361625 -96 -360649
rect -62 -361625 -50 -360649
rect -108 -361637 -50 -361625
rect 50 -360649 108 -360637
rect 50 -361625 62 -360649
rect 96 -361625 108 -360649
rect 50 -361637 108 -361625
rect -108 -361867 -50 -361855
rect -108 -362843 -96 -361867
rect -62 -362843 -50 -361867
rect -108 -362855 -50 -362843
rect 50 -361867 108 -361855
rect 50 -362843 62 -361867
rect 96 -362843 108 -361867
rect 50 -362855 108 -362843
rect -108 -363085 -50 -363073
rect -108 -364061 -96 -363085
rect -62 -364061 -50 -363085
rect -108 -364073 -50 -364061
rect 50 -363085 108 -363073
rect 50 -364061 62 -363085
rect 96 -364061 108 -363085
rect 50 -364073 108 -364061
rect -108 -364303 -50 -364291
rect -108 -365279 -96 -364303
rect -62 -365279 -50 -364303
rect -108 -365291 -50 -365279
rect 50 -364303 108 -364291
rect 50 -365279 62 -364303
rect 96 -365279 108 -364303
rect 50 -365291 108 -365279
rect -108 -365521 -50 -365509
rect -108 -366497 -96 -365521
rect -62 -366497 -50 -365521
rect -108 -366509 -50 -366497
rect 50 -365521 108 -365509
rect 50 -366497 62 -365521
rect 96 -366497 108 -365521
rect 50 -366509 108 -366497
rect -108 -366739 -50 -366727
rect -108 -367715 -96 -366739
rect -62 -367715 -50 -366739
rect -108 -367727 -50 -367715
rect 50 -366739 108 -366727
rect 50 -367715 62 -366739
rect 96 -367715 108 -366739
rect 50 -367727 108 -367715
rect -108 -367957 -50 -367945
rect -108 -368933 -96 -367957
rect -62 -368933 -50 -367957
rect -108 -368945 -50 -368933
rect 50 -367957 108 -367945
rect 50 -368933 62 -367957
rect 96 -368933 108 -367957
rect 50 -368945 108 -368933
rect -108 -369175 -50 -369163
rect -108 -370151 -96 -369175
rect -62 -370151 -50 -369175
rect -108 -370163 -50 -370151
rect 50 -369175 108 -369163
rect 50 -370151 62 -369175
rect 96 -370151 108 -369175
rect 50 -370163 108 -370151
rect -108 -370393 -50 -370381
rect -108 -371369 -96 -370393
rect -62 -371369 -50 -370393
rect -108 -371381 -50 -371369
rect 50 -370393 108 -370381
rect 50 -371369 62 -370393
rect 96 -371369 108 -370393
rect 50 -371381 108 -371369
rect -108 -371611 -50 -371599
rect -108 -372587 -96 -371611
rect -62 -372587 -50 -371611
rect -108 -372599 -50 -372587
rect 50 -371611 108 -371599
rect 50 -372587 62 -371611
rect 96 -372587 108 -371611
rect 50 -372599 108 -372587
rect -108 -372829 -50 -372817
rect -108 -373805 -96 -372829
rect -62 -373805 -50 -372829
rect -108 -373817 -50 -373805
rect 50 -372829 108 -372817
rect 50 -373805 62 -372829
rect 96 -373805 108 -372829
rect 50 -373817 108 -373805
rect -108 -374047 -50 -374035
rect -108 -375023 -96 -374047
rect -62 -375023 -50 -374047
rect -108 -375035 -50 -375023
rect 50 -374047 108 -374035
rect 50 -375023 62 -374047
rect 96 -375023 108 -374047
rect 50 -375035 108 -375023
rect -108 -375265 -50 -375253
rect -108 -376241 -96 -375265
rect -62 -376241 -50 -375265
rect -108 -376253 -50 -376241
rect 50 -375265 108 -375253
rect 50 -376241 62 -375265
rect 96 -376241 108 -375265
rect 50 -376253 108 -376241
rect -108 -376483 -50 -376471
rect -108 -377459 -96 -376483
rect -62 -377459 -50 -376483
rect -108 -377471 -50 -377459
rect 50 -376483 108 -376471
rect 50 -377459 62 -376483
rect 96 -377459 108 -376483
rect 50 -377471 108 -377459
rect -108 -377701 -50 -377689
rect -108 -378677 -96 -377701
rect -62 -378677 -50 -377701
rect -108 -378689 -50 -378677
rect 50 -377701 108 -377689
rect 50 -378677 62 -377701
rect 96 -378677 108 -377701
rect 50 -378689 108 -378677
rect -108 -378919 -50 -378907
rect -108 -379895 -96 -378919
rect -62 -379895 -50 -378919
rect -108 -379907 -50 -379895
rect 50 -378919 108 -378907
rect 50 -379895 62 -378919
rect 96 -379895 108 -378919
rect 50 -379907 108 -379895
rect -108 -380137 -50 -380125
rect -108 -381113 -96 -380137
rect -62 -381113 -50 -380137
rect -108 -381125 -50 -381113
rect 50 -380137 108 -380125
rect 50 -381113 62 -380137
rect 96 -381113 108 -380137
rect 50 -381125 108 -381113
rect -108 -381355 -50 -381343
rect -108 -382331 -96 -381355
rect -62 -382331 -50 -381355
rect -108 -382343 -50 -382331
rect 50 -381355 108 -381343
rect 50 -382331 62 -381355
rect 96 -382331 108 -381355
rect 50 -382343 108 -382331
rect -108 -382573 -50 -382561
rect -108 -383549 -96 -382573
rect -62 -383549 -50 -382573
rect -108 -383561 -50 -383549
rect 50 -382573 108 -382561
rect 50 -383549 62 -382573
rect 96 -383549 108 -382573
rect 50 -383561 108 -383549
rect -108 -383791 -50 -383779
rect -108 -384767 -96 -383791
rect -62 -384767 -50 -383791
rect -108 -384779 -50 -384767
rect 50 -383791 108 -383779
rect 50 -384767 62 -383791
rect 96 -384767 108 -383791
rect 50 -384779 108 -384767
rect -108 -385009 -50 -384997
rect -108 -385985 -96 -385009
rect -62 -385985 -50 -385009
rect -108 -385997 -50 -385985
rect 50 -385009 108 -384997
rect 50 -385985 62 -385009
rect 96 -385985 108 -385009
rect 50 -385997 108 -385985
rect -108 -386227 -50 -386215
rect -108 -387203 -96 -386227
rect -62 -387203 -50 -386227
rect -108 -387215 -50 -387203
rect 50 -386227 108 -386215
rect 50 -387203 62 -386227
rect 96 -387203 108 -386227
rect 50 -387215 108 -387203
rect -108 -387445 -50 -387433
rect -108 -388421 -96 -387445
rect -62 -388421 -50 -387445
rect -108 -388433 -50 -388421
rect 50 -387445 108 -387433
rect 50 -388421 62 -387445
rect 96 -388421 108 -387445
rect 50 -388433 108 -388421
rect -108 -388663 -50 -388651
rect -108 -389639 -96 -388663
rect -62 -389639 -50 -388663
rect -108 -389651 -50 -389639
rect 50 -388663 108 -388651
rect 50 -389639 62 -388663
rect 96 -389639 108 -388663
rect 50 -389651 108 -389639
rect -108 -389881 -50 -389869
rect -108 -390857 -96 -389881
rect -62 -390857 -50 -389881
rect -108 -390869 -50 -390857
rect 50 -389881 108 -389869
rect 50 -390857 62 -389881
rect 96 -390857 108 -389881
rect 50 -390869 108 -390857
rect -108 -391099 -50 -391087
rect -108 -392075 -96 -391099
rect -62 -392075 -50 -391099
rect -108 -392087 -50 -392075
rect 50 -391099 108 -391087
rect 50 -392075 62 -391099
rect 96 -392075 108 -391099
rect 50 -392087 108 -392075
rect -108 -392317 -50 -392305
rect -108 -393293 -96 -392317
rect -62 -393293 -50 -392317
rect -108 -393305 -50 -393293
rect 50 -392317 108 -392305
rect 50 -393293 62 -392317
rect 96 -393293 108 -392317
rect 50 -393305 108 -393293
rect -108 -393535 -50 -393523
rect -108 -394511 -96 -393535
rect -62 -394511 -50 -393535
rect -108 -394523 -50 -394511
rect 50 -393535 108 -393523
rect 50 -394511 62 -393535
rect 96 -394511 108 -393535
rect 50 -394523 108 -394511
rect -108 -394753 -50 -394741
rect -108 -395729 -96 -394753
rect -62 -395729 -50 -394753
rect -108 -395741 -50 -395729
rect 50 -394753 108 -394741
rect 50 -395729 62 -394753
rect 96 -395729 108 -394753
rect 50 -395741 108 -395729
rect -108 -395971 -50 -395959
rect -108 -396947 -96 -395971
rect -62 -396947 -50 -395971
rect -108 -396959 -50 -396947
rect 50 -395971 108 -395959
rect 50 -396947 62 -395971
rect 96 -396947 108 -395971
rect 50 -396959 108 -396947
rect -108 -397189 -50 -397177
rect -108 -398165 -96 -397189
rect -62 -398165 -50 -397189
rect -108 -398177 -50 -398165
rect 50 -397189 108 -397177
rect 50 -398165 62 -397189
rect 96 -398165 108 -397189
rect 50 -398177 108 -398165
rect -108 -398407 -50 -398395
rect -108 -399383 -96 -398407
rect -62 -399383 -50 -398407
rect -108 -399395 -50 -399383
rect 50 -398407 108 -398395
rect 50 -399383 62 -398407
rect 96 -399383 108 -398407
rect 50 -399395 108 -399383
rect -108 -399625 -50 -399613
rect -108 -400601 -96 -399625
rect -62 -400601 -50 -399625
rect -108 -400613 -50 -400601
rect 50 -399625 108 -399613
rect 50 -400601 62 -399625
rect 96 -400601 108 -399625
rect 50 -400613 108 -400601
rect -108 -400843 -50 -400831
rect -108 -401819 -96 -400843
rect -62 -401819 -50 -400843
rect -108 -401831 -50 -401819
rect 50 -400843 108 -400831
rect 50 -401819 62 -400843
rect 96 -401819 108 -400843
rect 50 -401831 108 -401819
rect -108 -402061 -50 -402049
rect -108 -403037 -96 -402061
rect -62 -403037 -50 -402061
rect -108 -403049 -50 -403037
rect 50 -402061 108 -402049
rect 50 -403037 62 -402061
rect 96 -403037 108 -402061
rect 50 -403049 108 -403037
rect -108 -403279 -50 -403267
rect -108 -404255 -96 -403279
rect -62 -404255 -50 -403279
rect -108 -404267 -50 -404255
rect 50 -403279 108 -403267
rect 50 -404255 62 -403279
rect 96 -404255 108 -403279
rect 50 -404267 108 -404255
rect -108 -404497 -50 -404485
rect -108 -405473 -96 -404497
rect -62 -405473 -50 -404497
rect -108 -405485 -50 -405473
rect 50 -404497 108 -404485
rect 50 -405473 62 -404497
rect 96 -405473 108 -404497
rect 50 -405485 108 -405473
rect -108 -405715 -50 -405703
rect -108 -406691 -96 -405715
rect -62 -406691 -50 -405715
rect -108 -406703 -50 -406691
rect 50 -405715 108 -405703
rect 50 -406691 62 -405715
rect 96 -406691 108 -405715
rect 50 -406703 108 -406691
rect -108 -406933 -50 -406921
rect -108 -407909 -96 -406933
rect -62 -407909 -50 -406933
rect -108 -407921 -50 -407909
rect 50 -406933 108 -406921
rect 50 -407909 62 -406933
rect 96 -407909 108 -406933
rect 50 -407921 108 -407909
rect -108 -408151 -50 -408139
rect -108 -409127 -96 -408151
rect -62 -409127 -50 -408151
rect -108 -409139 -50 -409127
rect 50 -408151 108 -408139
rect 50 -409127 62 -408151
rect 96 -409127 108 -408151
rect 50 -409139 108 -409127
rect -108 -409369 -50 -409357
rect -108 -410345 -96 -409369
rect -62 -410345 -50 -409369
rect -108 -410357 -50 -410345
rect 50 -409369 108 -409357
rect 50 -410345 62 -409369
rect 96 -410345 108 -409369
rect 50 -410357 108 -410345
rect -108 -410587 -50 -410575
rect -108 -411563 -96 -410587
rect -62 -411563 -50 -410587
rect -108 -411575 -50 -411563
rect 50 -410587 108 -410575
rect 50 -411563 62 -410587
rect 96 -411563 108 -410587
rect 50 -411575 108 -411563
rect -108 -411805 -50 -411793
rect -108 -412781 -96 -411805
rect -62 -412781 -50 -411805
rect -108 -412793 -50 -412781
rect 50 -411805 108 -411793
rect 50 -412781 62 -411805
rect 96 -412781 108 -411805
rect 50 -412793 108 -412781
rect -108 -413023 -50 -413011
rect -108 -413999 -96 -413023
rect -62 -413999 -50 -413023
rect -108 -414011 -50 -413999
rect 50 -413023 108 -413011
rect 50 -413999 62 -413023
rect 96 -413999 108 -413023
rect 50 -414011 108 -413999
rect -108 -414241 -50 -414229
rect -108 -415217 -96 -414241
rect -62 -415217 -50 -414241
rect -108 -415229 -50 -415217
rect 50 -414241 108 -414229
rect 50 -415217 62 -414241
rect 96 -415217 108 -414241
rect 50 -415229 108 -415217
rect -108 -415459 -50 -415447
rect -108 -416435 -96 -415459
rect -62 -416435 -50 -415459
rect -108 -416447 -50 -416435
rect 50 -415459 108 -415447
rect 50 -416435 62 -415459
rect 96 -416435 108 -415459
rect 50 -416447 108 -416435
rect -108 -416677 -50 -416665
rect -108 -417653 -96 -416677
rect -62 -417653 -50 -416677
rect -108 -417665 -50 -417653
rect 50 -416677 108 -416665
rect 50 -417653 62 -416677
rect 96 -417653 108 -416677
rect 50 -417665 108 -417653
rect -108 -417895 -50 -417883
rect -108 -418871 -96 -417895
rect -62 -418871 -50 -417895
rect -108 -418883 -50 -418871
rect 50 -417895 108 -417883
rect 50 -418871 62 -417895
rect 96 -418871 108 -417895
rect 50 -418883 108 -418871
rect -108 -419113 -50 -419101
rect -108 -420089 -96 -419113
rect -62 -420089 -50 -419113
rect -108 -420101 -50 -420089
rect 50 -419113 108 -419101
rect 50 -420089 62 -419113
rect 96 -420089 108 -419113
rect 50 -420101 108 -420089
rect -108 -420331 -50 -420319
rect -108 -421307 -96 -420331
rect -62 -421307 -50 -420331
rect -108 -421319 -50 -421307
rect 50 -420331 108 -420319
rect 50 -421307 62 -420331
rect 96 -421307 108 -420331
rect 50 -421319 108 -421307
rect -108 -421549 -50 -421537
rect -108 -422525 -96 -421549
rect -62 -422525 -50 -421549
rect -108 -422537 -50 -422525
rect 50 -421549 108 -421537
rect 50 -422525 62 -421549
rect 96 -422525 108 -421549
rect 50 -422537 108 -422525
rect -108 -422767 -50 -422755
rect -108 -423743 -96 -422767
rect -62 -423743 -50 -422767
rect -108 -423755 -50 -423743
rect 50 -422767 108 -422755
rect 50 -423743 62 -422767
rect 96 -423743 108 -422767
rect 50 -423755 108 -423743
rect -108 -423985 -50 -423973
rect -108 -424961 -96 -423985
rect -62 -424961 -50 -423985
rect -108 -424973 -50 -424961
rect 50 -423985 108 -423973
rect 50 -424961 62 -423985
rect 96 -424961 108 -423985
rect 50 -424973 108 -424961
rect -108 -425203 -50 -425191
rect -108 -426179 -96 -425203
rect -62 -426179 -50 -425203
rect -108 -426191 -50 -426179
rect 50 -425203 108 -425191
rect 50 -426179 62 -425203
rect 96 -426179 108 -425203
rect 50 -426191 108 -426179
rect -108 -426421 -50 -426409
rect -108 -427397 -96 -426421
rect -62 -427397 -50 -426421
rect -108 -427409 -50 -427397
rect 50 -426421 108 -426409
rect 50 -427397 62 -426421
rect 96 -427397 108 -426421
rect 50 -427409 108 -427397
rect -108 -427639 -50 -427627
rect -108 -428615 -96 -427639
rect -62 -428615 -50 -427639
rect -108 -428627 -50 -428615
rect 50 -427639 108 -427627
rect 50 -428615 62 -427639
rect 96 -428615 108 -427639
rect 50 -428627 108 -428615
rect -108 -428857 -50 -428845
rect -108 -429833 -96 -428857
rect -62 -429833 -50 -428857
rect -108 -429845 -50 -429833
rect 50 -428857 108 -428845
rect 50 -429833 62 -428857
rect 96 -429833 108 -428857
rect 50 -429845 108 -429833
rect -108 -430075 -50 -430063
rect -108 -431051 -96 -430075
rect -62 -431051 -50 -430075
rect -108 -431063 -50 -431051
rect 50 -430075 108 -430063
rect 50 -431051 62 -430075
rect 96 -431051 108 -430075
rect 50 -431063 108 -431051
rect -108 -431293 -50 -431281
rect -108 -432269 -96 -431293
rect -62 -432269 -50 -431293
rect -108 -432281 -50 -432269
rect 50 -431293 108 -431281
rect 50 -432269 62 -431293
rect 96 -432269 108 -431293
rect 50 -432281 108 -432269
rect -108 -432511 -50 -432499
rect -108 -433487 -96 -432511
rect -62 -433487 -50 -432511
rect -108 -433499 -50 -433487
rect 50 -432511 108 -432499
rect 50 -433487 62 -432511
rect 96 -433487 108 -432511
rect 50 -433499 108 -433487
rect -108 -433729 -50 -433717
rect -108 -434705 -96 -433729
rect -62 -434705 -50 -433729
rect -108 -434717 -50 -434705
rect 50 -433729 108 -433717
rect 50 -434705 62 -433729
rect 96 -434705 108 -433729
rect 50 -434717 108 -434705
rect -108 -434947 -50 -434935
rect -108 -435923 -96 -434947
rect -62 -435923 -50 -434947
rect -108 -435935 -50 -435923
rect 50 -434947 108 -434935
rect 50 -435923 62 -434947
rect 96 -435923 108 -434947
rect 50 -435935 108 -435923
rect -108 -436165 -50 -436153
rect -108 -437141 -96 -436165
rect -62 -437141 -50 -436165
rect -108 -437153 -50 -437141
rect 50 -436165 108 -436153
rect 50 -437141 62 -436165
rect 96 -437141 108 -436165
rect 50 -437153 108 -437141
rect -108 -437383 -50 -437371
rect -108 -438359 -96 -437383
rect -62 -438359 -50 -437383
rect -108 -438371 -50 -438359
rect 50 -437383 108 -437371
rect 50 -438359 62 -437383
rect 96 -438359 108 -437383
rect 50 -438371 108 -438359
rect -108 -438601 -50 -438589
rect -108 -439577 -96 -438601
rect -62 -439577 -50 -438601
rect -108 -439589 -50 -439577
rect 50 -438601 108 -438589
rect 50 -439577 62 -438601
rect 96 -439577 108 -438601
rect 50 -439589 108 -439577
rect -108 -439819 -50 -439807
rect -108 -440795 -96 -439819
rect -62 -440795 -50 -439819
rect -108 -440807 -50 -440795
rect 50 -439819 108 -439807
rect 50 -440795 62 -439819
rect 96 -440795 108 -439819
rect 50 -440807 108 -440795
rect -108 -441037 -50 -441025
rect -108 -442013 -96 -441037
rect -62 -442013 -50 -441037
rect -108 -442025 -50 -442013
rect 50 -441037 108 -441025
rect 50 -442013 62 -441037
rect 96 -442013 108 -441037
rect 50 -442025 108 -442013
rect -108 -442255 -50 -442243
rect -108 -443231 -96 -442255
rect -62 -443231 -50 -442255
rect -108 -443243 -50 -443231
rect 50 -442255 108 -442243
rect 50 -443231 62 -442255
rect 96 -443231 108 -442255
rect 50 -443243 108 -443231
rect -108 -443473 -50 -443461
rect -108 -444449 -96 -443473
rect -62 -444449 -50 -443473
rect -108 -444461 -50 -444449
rect 50 -443473 108 -443461
rect 50 -444449 62 -443473
rect 96 -444449 108 -443473
rect 50 -444461 108 -444449
rect -108 -444691 -50 -444679
rect -108 -445667 -96 -444691
rect -62 -445667 -50 -444691
rect -108 -445679 -50 -445667
rect 50 -444691 108 -444679
rect 50 -445667 62 -444691
rect 96 -445667 108 -444691
rect 50 -445679 108 -445667
rect -108 -445909 -50 -445897
rect -108 -446885 -96 -445909
rect -62 -446885 -50 -445909
rect -108 -446897 -50 -446885
rect 50 -445909 108 -445897
rect 50 -446885 62 -445909
rect 96 -446885 108 -445909
rect 50 -446897 108 -446885
rect -108 -447127 -50 -447115
rect -108 -448103 -96 -447127
rect -62 -448103 -50 -447127
rect -108 -448115 -50 -448103
rect 50 -447127 108 -447115
rect 50 -448103 62 -447127
rect 96 -448103 108 -447127
rect 50 -448115 108 -448103
rect -108 -448345 -50 -448333
rect -108 -449321 -96 -448345
rect -62 -449321 -50 -448345
rect -108 -449333 -50 -449321
rect 50 -448345 108 -448333
rect 50 -449321 62 -448345
rect 96 -449321 108 -448345
rect 50 -449333 108 -449321
rect -108 -449563 -50 -449551
rect -108 -450539 -96 -449563
rect -62 -450539 -50 -449563
rect -108 -450551 -50 -450539
rect 50 -449563 108 -449551
rect 50 -450539 62 -449563
rect 96 -450539 108 -449563
rect 50 -450551 108 -450539
rect -108 -450781 -50 -450769
rect -108 -451757 -96 -450781
rect -62 -451757 -50 -450781
rect -108 -451769 -50 -451757
rect 50 -450781 108 -450769
rect 50 -451757 62 -450781
rect 96 -451757 108 -450781
rect 50 -451769 108 -451757
rect -108 -451999 -50 -451987
rect -108 -452975 -96 -451999
rect -62 -452975 -50 -451999
rect -108 -452987 -50 -452975
rect 50 -451999 108 -451987
rect 50 -452975 62 -451999
rect 96 -452975 108 -451999
rect 50 -452987 108 -452975
rect -108 -453217 -50 -453205
rect -108 -454193 -96 -453217
rect -62 -454193 -50 -453217
rect -108 -454205 -50 -454193
rect 50 -453217 108 -453205
rect 50 -454193 62 -453217
rect 96 -454193 108 -453217
rect 50 -454205 108 -454193
rect -108 -454435 -50 -454423
rect -108 -455411 -96 -454435
rect -62 -455411 -50 -454435
rect -108 -455423 -50 -455411
rect 50 -454435 108 -454423
rect 50 -455411 62 -454435
rect 96 -455411 108 -454435
rect 50 -455423 108 -455411
rect -108 -455653 -50 -455641
rect -108 -456629 -96 -455653
rect -62 -456629 -50 -455653
rect -108 -456641 -50 -456629
rect 50 -455653 108 -455641
rect 50 -456629 62 -455653
rect 96 -456629 108 -455653
rect 50 -456641 108 -456629
rect -108 -456871 -50 -456859
rect -108 -457847 -96 -456871
rect -62 -457847 -50 -456871
rect -108 -457859 -50 -457847
rect 50 -456871 108 -456859
rect 50 -457847 62 -456871
rect 96 -457847 108 -456871
rect 50 -457859 108 -457847
rect -108 -458089 -50 -458077
rect -108 -459065 -96 -458089
rect -62 -459065 -50 -458089
rect -108 -459077 -50 -459065
rect 50 -458089 108 -458077
rect 50 -459065 62 -458089
rect 96 -459065 108 -458089
rect 50 -459077 108 -459065
rect -108 -459307 -50 -459295
rect -108 -460283 -96 -459307
rect -62 -460283 -50 -459307
rect -108 -460295 -50 -460283
rect 50 -459307 108 -459295
rect 50 -460283 62 -459307
rect 96 -460283 108 -459307
rect 50 -460295 108 -460283
rect -108 -460525 -50 -460513
rect -108 -461501 -96 -460525
rect -62 -461501 -50 -460525
rect -108 -461513 -50 -461501
rect 50 -460525 108 -460513
rect 50 -461501 62 -460525
rect 96 -461501 108 -460525
rect 50 -461513 108 -461501
rect -108 -461743 -50 -461731
rect -108 -462719 -96 -461743
rect -62 -462719 -50 -461743
rect -108 -462731 -50 -462719
rect 50 -461743 108 -461731
rect 50 -462719 62 -461743
rect 96 -462719 108 -461743
rect 50 -462731 108 -462719
rect -108 -462961 -50 -462949
rect -108 -463937 -96 -462961
rect -62 -463937 -50 -462961
rect -108 -463949 -50 -463937
rect 50 -462961 108 -462949
rect 50 -463937 62 -462961
rect 96 -463937 108 -462961
rect 50 -463949 108 -463937
rect -108 -464179 -50 -464167
rect -108 -465155 -96 -464179
rect -62 -465155 -50 -464179
rect -108 -465167 -50 -465155
rect 50 -464179 108 -464167
rect 50 -465155 62 -464179
rect 96 -465155 108 -464179
rect 50 -465167 108 -465155
rect -108 -465397 -50 -465385
rect -108 -466373 -96 -465397
rect -62 -466373 -50 -465397
rect -108 -466385 -50 -466373
rect 50 -465397 108 -465385
rect 50 -466373 62 -465397
rect 96 -466373 108 -465397
rect 50 -466385 108 -466373
rect -108 -466615 -50 -466603
rect -108 -467591 -96 -466615
rect -62 -467591 -50 -466615
rect -108 -467603 -50 -467591
rect 50 -466615 108 -466603
rect 50 -467591 62 -466615
rect 96 -467591 108 -466615
rect 50 -467603 108 -467591
rect -108 -467833 -50 -467821
rect -108 -468809 -96 -467833
rect -62 -468809 -50 -467833
rect -108 -468821 -50 -468809
rect 50 -467833 108 -467821
rect 50 -468809 62 -467833
rect 96 -468809 108 -467833
rect 50 -468821 108 -468809
rect -108 -469051 -50 -469039
rect -108 -470027 -96 -469051
rect -62 -470027 -50 -469051
rect -108 -470039 -50 -470027
rect 50 -469051 108 -469039
rect 50 -470027 62 -469051
rect 96 -470027 108 -469051
rect 50 -470039 108 -470027
rect -108 -470269 -50 -470257
rect -108 -471245 -96 -470269
rect -62 -471245 -50 -470269
rect -108 -471257 -50 -471245
rect 50 -470269 108 -470257
rect 50 -471245 62 -470269
rect 96 -471245 108 -470269
rect 50 -471257 108 -471245
rect -108 -471487 -50 -471475
rect -108 -472463 -96 -471487
rect -62 -472463 -50 -471487
rect -108 -472475 -50 -472463
rect 50 -471487 108 -471475
rect 50 -472463 62 -471487
rect 96 -472463 108 -471487
rect 50 -472475 108 -472463
rect -108 -472705 -50 -472693
rect -108 -473681 -96 -472705
rect -62 -473681 -50 -472705
rect -108 -473693 -50 -473681
rect 50 -472705 108 -472693
rect 50 -473681 62 -472705
rect 96 -473681 108 -472705
rect 50 -473693 108 -473681
rect -108 -473923 -50 -473911
rect -108 -474899 -96 -473923
rect -62 -474899 -50 -473923
rect -108 -474911 -50 -474899
rect 50 -473923 108 -473911
rect 50 -474899 62 -473923
rect 96 -474899 108 -473923
rect 50 -474911 108 -474899
rect -108 -475141 -50 -475129
rect -108 -476117 -96 -475141
rect -62 -476117 -50 -475141
rect -108 -476129 -50 -476117
rect 50 -475141 108 -475129
rect 50 -476117 62 -475141
rect 96 -476117 108 -475141
rect 50 -476129 108 -476117
rect -108 -476359 -50 -476347
rect -108 -477335 -96 -476359
rect -62 -477335 -50 -476359
rect -108 -477347 -50 -477335
rect 50 -476359 108 -476347
rect 50 -477335 62 -476359
rect 96 -477335 108 -476359
rect 50 -477347 108 -477335
rect -108 -477577 -50 -477565
rect -108 -478553 -96 -477577
rect -62 -478553 -50 -477577
rect -108 -478565 -50 -478553
rect 50 -477577 108 -477565
rect 50 -478553 62 -477577
rect 96 -478553 108 -477577
rect 50 -478565 108 -478553
rect -108 -478795 -50 -478783
rect -108 -479771 -96 -478795
rect -62 -479771 -50 -478795
rect -108 -479783 -50 -479771
rect 50 -478795 108 -478783
rect 50 -479771 62 -478795
rect 96 -479771 108 -478795
rect 50 -479783 108 -479771
rect -108 -480013 -50 -480001
rect -108 -480989 -96 -480013
rect -62 -480989 -50 -480013
rect -108 -481001 -50 -480989
rect 50 -480013 108 -480001
rect 50 -480989 62 -480013
rect 96 -480989 108 -480013
rect 50 -481001 108 -480989
rect -108 -481231 -50 -481219
rect -108 -482207 -96 -481231
rect -62 -482207 -50 -481231
rect -108 -482219 -50 -482207
rect 50 -481231 108 -481219
rect 50 -482207 62 -481231
rect 96 -482207 108 -481231
rect 50 -482219 108 -482207
rect -108 -482449 -50 -482437
rect -108 -483425 -96 -482449
rect -62 -483425 -50 -482449
rect -108 -483437 -50 -483425
rect 50 -482449 108 -482437
rect 50 -483425 62 -482449
rect 96 -483425 108 -482449
rect 50 -483437 108 -483425
rect -108 -483667 -50 -483655
rect -108 -484643 -96 -483667
rect -62 -484643 -50 -483667
rect -108 -484655 -50 -484643
rect 50 -483667 108 -483655
rect 50 -484643 62 -483667
rect 96 -484643 108 -483667
rect 50 -484655 108 -484643
rect -108 -484885 -50 -484873
rect -108 -485861 -96 -484885
rect -62 -485861 -50 -484885
rect -108 -485873 -50 -485861
rect 50 -484885 108 -484873
rect 50 -485861 62 -484885
rect 96 -485861 108 -484885
rect 50 -485873 108 -485861
rect -108 -486103 -50 -486091
rect -108 -487079 -96 -486103
rect -62 -487079 -50 -486103
rect -108 -487091 -50 -487079
rect 50 -486103 108 -486091
rect 50 -487079 62 -486103
rect 96 -487079 108 -486103
rect 50 -487091 108 -487079
rect -108 -487321 -50 -487309
rect -108 -488297 -96 -487321
rect -62 -488297 -50 -487321
rect -108 -488309 -50 -488297
rect 50 -487321 108 -487309
rect 50 -488297 62 -487321
rect 96 -488297 108 -487321
rect 50 -488309 108 -488297
rect -108 -488539 -50 -488527
rect -108 -489515 -96 -488539
rect -62 -489515 -50 -488539
rect -108 -489527 -50 -489515
rect 50 -488539 108 -488527
rect 50 -489515 62 -488539
rect 96 -489515 108 -488539
rect 50 -489527 108 -489515
rect -108 -489757 -50 -489745
rect -108 -490733 -96 -489757
rect -62 -490733 -50 -489757
rect -108 -490745 -50 -490733
rect 50 -489757 108 -489745
rect 50 -490733 62 -489757
rect 96 -490733 108 -489757
rect 50 -490745 108 -490733
rect -108 -490975 -50 -490963
rect -108 -491951 -96 -490975
rect -62 -491951 -50 -490975
rect -108 -491963 -50 -491951
rect 50 -490975 108 -490963
rect 50 -491951 62 -490975
rect 96 -491951 108 -490975
rect 50 -491963 108 -491951
rect -108 -492193 -50 -492181
rect -108 -493169 -96 -492193
rect -62 -493169 -50 -492193
rect -108 -493181 -50 -493169
rect 50 -492193 108 -492181
rect 50 -493169 62 -492193
rect 96 -493169 108 -492193
rect 50 -493181 108 -493169
rect -108 -493411 -50 -493399
rect -108 -494387 -96 -493411
rect -62 -494387 -50 -493411
rect -108 -494399 -50 -494387
rect 50 -493411 108 -493399
rect 50 -494387 62 -493411
rect 96 -494387 108 -493411
rect 50 -494399 108 -494387
rect -108 -494629 -50 -494617
rect -108 -495605 -96 -494629
rect -62 -495605 -50 -494629
rect -108 -495617 -50 -495605
rect 50 -494629 108 -494617
rect 50 -495605 62 -494629
rect 96 -495605 108 -494629
rect 50 -495617 108 -495605
rect -108 -495847 -50 -495835
rect -108 -496823 -96 -495847
rect -62 -496823 -50 -495847
rect -108 -496835 -50 -496823
rect 50 -495847 108 -495835
rect 50 -496823 62 -495847
rect 96 -496823 108 -495847
rect 50 -496835 108 -496823
rect -108 -497065 -50 -497053
rect -108 -498041 -96 -497065
rect -62 -498041 -50 -497065
rect -108 -498053 -50 -498041
rect 50 -497065 108 -497053
rect 50 -498041 62 -497065
rect 96 -498041 108 -497065
rect 50 -498053 108 -498041
rect -108 -498283 -50 -498271
rect -108 -499259 -96 -498283
rect -62 -499259 -50 -498283
rect -108 -499271 -50 -499259
rect 50 -498283 108 -498271
rect 50 -499259 62 -498283
rect 96 -499259 108 -498283
rect 50 -499271 108 -499259
rect -108 -499501 -50 -499489
rect -108 -500477 -96 -499501
rect -62 -500477 -50 -499501
rect -108 -500489 -50 -500477
rect 50 -499501 108 -499489
rect 50 -500477 62 -499501
rect 96 -500477 108 -499501
rect 50 -500489 108 -500477
rect -108 -500719 -50 -500707
rect -108 -501695 -96 -500719
rect -62 -501695 -50 -500719
rect -108 -501707 -50 -501695
rect 50 -500719 108 -500707
rect 50 -501695 62 -500719
rect 96 -501695 108 -500719
rect 50 -501707 108 -501695
rect -108 -501937 -50 -501925
rect -108 -502913 -96 -501937
rect -62 -502913 -50 -501937
rect -108 -502925 -50 -502913
rect 50 -501937 108 -501925
rect 50 -502913 62 -501937
rect 96 -502913 108 -501937
rect 50 -502925 108 -502913
rect -108 -503155 -50 -503143
rect -108 -504131 -96 -503155
rect -62 -504131 -50 -503155
rect -108 -504143 -50 -504131
rect 50 -503155 108 -503143
rect 50 -504131 62 -503155
rect 96 -504131 108 -503155
rect 50 -504143 108 -504131
rect -108 -504373 -50 -504361
rect -108 -505349 -96 -504373
rect -62 -505349 -50 -504373
rect -108 -505361 -50 -505349
rect 50 -504373 108 -504361
rect 50 -505349 62 -504373
rect 96 -505349 108 -504373
rect 50 -505361 108 -505349
rect -108 -505591 -50 -505579
rect -108 -506567 -96 -505591
rect -62 -506567 -50 -505591
rect -108 -506579 -50 -506567
rect 50 -505591 108 -505579
rect 50 -506567 62 -505591
rect 96 -506567 108 -505591
rect 50 -506579 108 -506567
rect -108 -506809 -50 -506797
rect -108 -507785 -96 -506809
rect -62 -507785 -50 -506809
rect -108 -507797 -50 -507785
rect 50 -506809 108 -506797
rect 50 -507785 62 -506809
rect 96 -507785 108 -506809
rect 50 -507797 108 -507785
rect -108 -508027 -50 -508015
rect -108 -509003 -96 -508027
rect -62 -509003 -50 -508027
rect -108 -509015 -50 -509003
rect 50 -508027 108 -508015
rect 50 -509003 62 -508027
rect 96 -509003 108 -508027
rect 50 -509015 108 -509003
rect -108 -509245 -50 -509233
rect -108 -510221 -96 -509245
rect -62 -510221 -50 -509245
rect -108 -510233 -50 -510221
rect 50 -509245 108 -509233
rect 50 -510221 62 -509245
rect 96 -510221 108 -509245
rect 50 -510233 108 -510221
rect -108 -510463 -50 -510451
rect -108 -511439 -96 -510463
rect -62 -511439 -50 -510463
rect -108 -511451 -50 -511439
rect 50 -510463 108 -510451
rect 50 -511439 62 -510463
rect 96 -511439 108 -510463
rect 50 -511451 108 -511439
rect -108 -511681 -50 -511669
rect -108 -512657 -96 -511681
rect -62 -512657 -50 -511681
rect -108 -512669 -50 -512657
rect 50 -511681 108 -511669
rect 50 -512657 62 -511681
rect 96 -512657 108 -511681
rect 50 -512669 108 -512657
rect -108 -512899 -50 -512887
rect -108 -513875 -96 -512899
rect -62 -513875 -50 -512899
rect -108 -513887 -50 -513875
rect 50 -512899 108 -512887
rect 50 -513875 62 -512899
rect 96 -513875 108 -512899
rect 50 -513887 108 -513875
rect -108 -514117 -50 -514105
rect -108 -515093 -96 -514117
rect -62 -515093 -50 -514117
rect -108 -515105 -50 -515093
rect 50 -514117 108 -514105
rect 50 -515093 62 -514117
rect 96 -515093 108 -514117
rect 50 -515105 108 -515093
rect -108 -515335 -50 -515323
rect -108 -516311 -96 -515335
rect -62 -516311 -50 -515335
rect -108 -516323 -50 -516311
rect 50 -515335 108 -515323
rect 50 -516311 62 -515335
rect 96 -516311 108 -515335
rect 50 -516323 108 -516311
rect -108 -516553 -50 -516541
rect -108 -517529 -96 -516553
rect -62 -517529 -50 -516553
rect -108 -517541 -50 -517529
rect 50 -516553 108 -516541
rect 50 -517529 62 -516553
rect 96 -517529 108 -516553
rect 50 -517541 108 -517529
rect -108 -517771 -50 -517759
rect -108 -518747 -96 -517771
rect -62 -518747 -50 -517771
rect -108 -518759 -50 -518747
rect 50 -517771 108 -517759
rect 50 -518747 62 -517771
rect 96 -518747 108 -517771
rect 50 -518759 108 -518747
rect -108 -518989 -50 -518977
rect -108 -519965 -96 -518989
rect -62 -519965 -50 -518989
rect -108 -519977 -50 -519965
rect 50 -518989 108 -518977
rect 50 -519965 62 -518989
rect 96 -519965 108 -518989
rect 50 -519977 108 -519965
rect -108 -520207 -50 -520195
rect -108 -521183 -96 -520207
rect -62 -521183 -50 -520207
rect -108 -521195 -50 -521183
rect 50 -520207 108 -520195
rect 50 -521183 62 -520207
rect 96 -521183 108 -520207
rect 50 -521195 108 -521183
rect -108 -521425 -50 -521413
rect -108 -522401 -96 -521425
rect -62 -522401 -50 -521425
rect -108 -522413 -50 -522401
rect 50 -521425 108 -521413
rect 50 -522401 62 -521425
rect 96 -522401 108 -521425
rect 50 -522413 108 -522401
rect -108 -522643 -50 -522631
rect -108 -523619 -96 -522643
rect -62 -523619 -50 -522643
rect -108 -523631 -50 -523619
rect 50 -522643 108 -522631
rect 50 -523619 62 -522643
rect 96 -523619 108 -522643
rect 50 -523631 108 -523619
rect -108 -523861 -50 -523849
rect -108 -524837 -96 -523861
rect -62 -524837 -50 -523861
rect -108 -524849 -50 -524837
rect 50 -523861 108 -523849
rect 50 -524837 62 -523861
rect 96 -524837 108 -523861
rect 50 -524849 108 -524837
rect -108 -525079 -50 -525067
rect -108 -526055 -96 -525079
rect -62 -526055 -50 -525079
rect -108 -526067 -50 -526055
rect 50 -525079 108 -525067
rect 50 -526055 62 -525079
rect 96 -526055 108 -525079
rect 50 -526067 108 -526055
rect -108 -526297 -50 -526285
rect -108 -527273 -96 -526297
rect -62 -527273 -50 -526297
rect -108 -527285 -50 -527273
rect 50 -526297 108 -526285
rect 50 -527273 62 -526297
rect 96 -527273 108 -526297
rect 50 -527285 108 -527273
rect -108 -527515 -50 -527503
rect -108 -528491 -96 -527515
rect -62 -528491 -50 -527515
rect -108 -528503 -50 -528491
rect 50 -527515 108 -527503
rect 50 -528491 62 -527515
rect 96 -528491 108 -527515
rect 50 -528503 108 -528491
rect -108 -528733 -50 -528721
rect -108 -529709 -96 -528733
rect -62 -529709 -50 -528733
rect -108 -529721 -50 -529709
rect 50 -528733 108 -528721
rect 50 -529709 62 -528733
rect 96 -529709 108 -528733
rect 50 -529721 108 -529709
rect -108 -529951 -50 -529939
rect -108 -530927 -96 -529951
rect -62 -530927 -50 -529951
rect -108 -530939 -50 -530927
rect 50 -529951 108 -529939
rect 50 -530927 62 -529951
rect 96 -530927 108 -529951
rect 50 -530939 108 -530927
rect -108 -531169 -50 -531157
rect -108 -532145 -96 -531169
rect -62 -532145 -50 -531169
rect -108 -532157 -50 -532145
rect 50 -531169 108 -531157
rect 50 -532145 62 -531169
rect 96 -532145 108 -531169
rect 50 -532157 108 -532145
rect -108 -532387 -50 -532375
rect -108 -533363 -96 -532387
rect -62 -533363 -50 -532387
rect -108 -533375 -50 -533363
rect 50 -532387 108 -532375
rect 50 -533363 62 -532387
rect 96 -533363 108 -532387
rect 50 -533375 108 -533363
rect -108 -533605 -50 -533593
rect -108 -534581 -96 -533605
rect -62 -534581 -50 -533605
rect -108 -534593 -50 -534581
rect 50 -533605 108 -533593
rect 50 -534581 62 -533605
rect 96 -534581 108 -533605
rect 50 -534593 108 -534581
rect -108 -534823 -50 -534811
rect -108 -535799 -96 -534823
rect -62 -535799 -50 -534823
rect -108 -535811 -50 -535799
rect 50 -534823 108 -534811
rect 50 -535799 62 -534823
rect 96 -535799 108 -534823
rect 50 -535811 108 -535799
rect -108 -536041 -50 -536029
rect -108 -537017 -96 -536041
rect -62 -537017 -50 -536041
rect -108 -537029 -50 -537017
rect 50 -536041 108 -536029
rect 50 -537017 62 -536041
rect 96 -537017 108 -536041
rect 50 -537029 108 -537017
rect -108 -537259 -50 -537247
rect -108 -538235 -96 -537259
rect -62 -538235 -50 -537259
rect -108 -538247 -50 -538235
rect 50 -537259 108 -537247
rect 50 -538235 62 -537259
rect 96 -538235 108 -537259
rect 50 -538247 108 -538235
rect -108 -538477 -50 -538465
rect -108 -539453 -96 -538477
rect -62 -539453 -50 -538477
rect -108 -539465 -50 -539453
rect 50 -538477 108 -538465
rect 50 -539453 62 -538477
rect 96 -539453 108 -538477
rect 50 -539465 108 -539453
rect -108 -539695 -50 -539683
rect -108 -540671 -96 -539695
rect -62 -540671 -50 -539695
rect -108 -540683 -50 -540671
rect 50 -539695 108 -539683
rect 50 -540671 62 -539695
rect 96 -540671 108 -539695
rect 50 -540683 108 -540671
rect -108 -540913 -50 -540901
rect -108 -541889 -96 -540913
rect -62 -541889 -50 -540913
rect -108 -541901 -50 -541889
rect 50 -540913 108 -540901
rect 50 -541889 62 -540913
rect 96 -541889 108 -540913
rect 50 -541901 108 -541889
rect -108 -542131 -50 -542119
rect -108 -543107 -96 -542131
rect -62 -543107 -50 -542131
rect -108 -543119 -50 -543107
rect 50 -542131 108 -542119
rect 50 -543107 62 -542131
rect 96 -543107 108 -542131
rect 50 -543119 108 -543107
rect -108 -543349 -50 -543337
rect -108 -544325 -96 -543349
rect -62 -544325 -50 -543349
rect -108 -544337 -50 -544325
rect 50 -543349 108 -543337
rect 50 -544325 62 -543349
rect 96 -544325 108 -543349
rect 50 -544337 108 -544325
rect -108 -544567 -50 -544555
rect -108 -545543 -96 -544567
rect -62 -545543 -50 -544567
rect -108 -545555 -50 -545543
rect 50 -544567 108 -544555
rect 50 -545543 62 -544567
rect 96 -545543 108 -544567
rect 50 -545555 108 -545543
rect -108 -545785 -50 -545773
rect -108 -546761 -96 -545785
rect -62 -546761 -50 -545785
rect -108 -546773 -50 -546761
rect 50 -545785 108 -545773
rect 50 -546761 62 -545785
rect 96 -546761 108 -545785
rect 50 -546773 108 -546761
rect -108 -547003 -50 -546991
rect -108 -547979 -96 -547003
rect -62 -547979 -50 -547003
rect -108 -547991 -50 -547979
rect 50 -547003 108 -546991
rect 50 -547979 62 -547003
rect 96 -547979 108 -547003
rect 50 -547991 108 -547979
rect -108 -548221 -50 -548209
rect -108 -549197 -96 -548221
rect -62 -549197 -50 -548221
rect -108 -549209 -50 -549197
rect 50 -548221 108 -548209
rect 50 -549197 62 -548221
rect 96 -549197 108 -548221
rect 50 -549209 108 -549197
rect -108 -549439 -50 -549427
rect -108 -550415 -96 -549439
rect -62 -550415 -50 -549439
rect -108 -550427 -50 -550415
rect 50 -549439 108 -549427
rect 50 -550415 62 -549439
rect 96 -550415 108 -549439
rect 50 -550427 108 -550415
rect -108 -550657 -50 -550645
rect -108 -551633 -96 -550657
rect -62 -551633 -50 -550657
rect -108 -551645 -50 -551633
rect 50 -550657 108 -550645
rect 50 -551633 62 -550657
rect 96 -551633 108 -550657
rect 50 -551645 108 -551633
rect -108 -551875 -50 -551863
rect -108 -552851 -96 -551875
rect -62 -552851 -50 -551875
rect -108 -552863 -50 -552851
rect 50 -551875 108 -551863
rect 50 -552851 62 -551875
rect 96 -552851 108 -551875
rect 50 -552863 108 -552851
rect -108 -553093 -50 -553081
rect -108 -554069 -96 -553093
rect -62 -554069 -50 -553093
rect -108 -554081 -50 -554069
rect 50 -553093 108 -553081
rect 50 -554069 62 -553093
rect 96 -554069 108 -553093
rect 50 -554081 108 -554069
rect -108 -554311 -50 -554299
rect -108 -555287 -96 -554311
rect -62 -555287 -50 -554311
rect -108 -555299 -50 -555287
rect 50 -554311 108 -554299
rect 50 -555287 62 -554311
rect 96 -555287 108 -554311
rect 50 -555299 108 -555287
rect -108 -555529 -50 -555517
rect -108 -556505 -96 -555529
rect -62 -556505 -50 -555529
rect -108 -556517 -50 -556505
rect 50 -555529 108 -555517
rect 50 -556505 62 -555529
rect 96 -556505 108 -555529
rect 50 -556517 108 -556505
rect -108 -556747 -50 -556735
rect -108 -557723 -96 -556747
rect -62 -557723 -50 -556747
rect -108 -557735 -50 -557723
rect 50 -556747 108 -556735
rect 50 -557723 62 -556747
rect 96 -557723 108 -556747
rect 50 -557735 108 -557723
rect -108 -557965 -50 -557953
rect -108 -558941 -96 -557965
rect -62 -558941 -50 -557965
rect -108 -558953 -50 -558941
rect 50 -557965 108 -557953
rect 50 -558941 62 -557965
rect 96 -558941 108 -557965
rect 50 -558953 108 -558941
rect -108 -559183 -50 -559171
rect -108 -560159 -96 -559183
rect -62 -560159 -50 -559183
rect -108 -560171 -50 -560159
rect 50 -559183 108 -559171
rect 50 -560159 62 -559183
rect 96 -560159 108 -559183
rect 50 -560171 108 -560159
rect -108 -560401 -50 -560389
rect -108 -561377 -96 -560401
rect -62 -561377 -50 -560401
rect -108 -561389 -50 -561377
rect 50 -560401 108 -560389
rect 50 -561377 62 -560401
rect 96 -561377 108 -560401
rect 50 -561389 108 -561377
rect -108 -561619 -50 -561607
rect -108 -562595 -96 -561619
rect -62 -562595 -50 -561619
rect -108 -562607 -50 -562595
rect 50 -561619 108 -561607
rect 50 -562595 62 -561619
rect 96 -562595 108 -561619
rect 50 -562607 108 -562595
rect -108 -562837 -50 -562825
rect -108 -563813 -96 -562837
rect -62 -563813 -50 -562837
rect -108 -563825 -50 -563813
rect 50 -562837 108 -562825
rect 50 -563813 62 -562837
rect 96 -563813 108 -562837
rect 50 -563825 108 -563813
rect -108 -564055 -50 -564043
rect -108 -565031 -96 -564055
rect -62 -565031 -50 -564055
rect -108 -565043 -50 -565031
rect 50 -564055 108 -564043
rect 50 -565031 62 -564055
rect 96 -565031 108 -564055
rect 50 -565043 108 -565031
rect -108 -565273 -50 -565261
rect -108 -566249 -96 -565273
rect -62 -566249 -50 -565273
rect -108 -566261 -50 -566249
rect 50 -565273 108 -565261
rect 50 -566249 62 -565273
rect 96 -566249 108 -565273
rect 50 -566261 108 -566249
rect -108 -566491 -50 -566479
rect -108 -567467 -96 -566491
rect -62 -567467 -50 -566491
rect -108 -567479 -50 -567467
rect 50 -566491 108 -566479
rect 50 -567467 62 -566491
rect 96 -567467 108 -566491
rect 50 -567479 108 -567467
rect -108 -567709 -50 -567697
rect -108 -568685 -96 -567709
rect -62 -568685 -50 -567709
rect -108 -568697 -50 -568685
rect 50 -567709 108 -567697
rect 50 -568685 62 -567709
rect 96 -568685 108 -567709
rect 50 -568697 108 -568685
rect -108 -568927 -50 -568915
rect -108 -569903 -96 -568927
rect -62 -569903 -50 -568927
rect -108 -569915 -50 -569903
rect 50 -568927 108 -568915
rect 50 -569903 62 -568927
rect 96 -569903 108 -568927
rect 50 -569915 108 -569903
rect -108 -570145 -50 -570133
rect -108 -571121 -96 -570145
rect -62 -571121 -50 -570145
rect -108 -571133 -50 -571121
rect 50 -570145 108 -570133
rect 50 -571121 62 -570145
rect 96 -571121 108 -570145
rect 50 -571133 108 -571121
rect -108 -571363 -50 -571351
rect -108 -572339 -96 -571363
rect -62 -572339 -50 -571363
rect -108 -572351 -50 -572339
rect 50 -571363 108 -571351
rect 50 -572339 62 -571363
rect 96 -572339 108 -571363
rect 50 -572351 108 -572339
rect -108 -572581 -50 -572569
rect -108 -573557 -96 -572581
rect -62 -573557 -50 -572581
rect -108 -573569 -50 -573557
rect 50 -572581 108 -572569
rect 50 -573557 62 -572581
rect 96 -573557 108 -572581
rect 50 -573569 108 -573557
rect -108 -573799 -50 -573787
rect -108 -574775 -96 -573799
rect -62 -574775 -50 -573799
rect -108 -574787 -50 -574775
rect 50 -573799 108 -573787
rect 50 -574775 62 -573799
rect 96 -574775 108 -573799
rect 50 -574787 108 -574775
rect -108 -575017 -50 -575005
rect -108 -575993 -96 -575017
rect -62 -575993 -50 -575017
rect -108 -576005 -50 -575993
rect 50 -575017 108 -575005
rect 50 -575993 62 -575017
rect 96 -575993 108 -575017
rect 50 -576005 108 -575993
rect -108 -576235 -50 -576223
rect -108 -577211 -96 -576235
rect -62 -577211 -50 -576235
rect -108 -577223 -50 -577211
rect 50 -576235 108 -576223
rect 50 -577211 62 -576235
rect 96 -577211 108 -576235
rect 50 -577223 108 -577211
rect -108 -577453 -50 -577441
rect -108 -578429 -96 -577453
rect -62 -578429 -50 -577453
rect -108 -578441 -50 -578429
rect 50 -577453 108 -577441
rect 50 -578429 62 -577453
rect 96 -578429 108 -577453
rect 50 -578441 108 -578429
rect -108 -578671 -50 -578659
rect -108 -579647 -96 -578671
rect -62 -579647 -50 -578671
rect -108 -579659 -50 -579647
rect 50 -578671 108 -578659
rect 50 -579647 62 -578671
rect 96 -579647 108 -578671
rect 50 -579659 108 -579647
rect -108 -579889 -50 -579877
rect -108 -580865 -96 -579889
rect -62 -580865 -50 -579889
rect -108 -580877 -50 -580865
rect 50 -579889 108 -579877
rect 50 -580865 62 -579889
rect 96 -580865 108 -579889
rect 50 -580877 108 -580865
rect -108 -581107 -50 -581095
rect -108 -582083 -96 -581107
rect -62 -582083 -50 -581107
rect -108 -582095 -50 -582083
rect 50 -581107 108 -581095
rect 50 -582083 62 -581107
rect 96 -582083 108 -581107
rect 50 -582095 108 -582083
rect -108 -582325 -50 -582313
rect -108 -583301 -96 -582325
rect -62 -583301 -50 -582325
rect -108 -583313 -50 -583301
rect 50 -582325 108 -582313
rect 50 -583301 62 -582325
rect 96 -583301 108 -582325
rect 50 -583313 108 -583301
rect -108 -583543 -50 -583531
rect -108 -584519 -96 -583543
rect -62 -584519 -50 -583543
rect -108 -584531 -50 -584519
rect 50 -583543 108 -583531
rect 50 -584519 62 -583543
rect 96 -584519 108 -583543
rect 50 -584531 108 -584519
rect -108 -584761 -50 -584749
rect -108 -585737 -96 -584761
rect -62 -585737 -50 -584761
rect -108 -585749 -50 -585737
rect 50 -584761 108 -584749
rect 50 -585737 62 -584761
rect 96 -585737 108 -584761
rect 50 -585749 108 -585737
rect -108 -585979 -50 -585967
rect -108 -586955 -96 -585979
rect -62 -586955 -50 -585979
rect -108 -586967 -50 -586955
rect 50 -585979 108 -585967
rect 50 -586955 62 -585979
rect 96 -586955 108 -585979
rect 50 -586967 108 -586955
rect -108 -587197 -50 -587185
rect -108 -588173 -96 -587197
rect -62 -588173 -50 -587197
rect -108 -588185 -50 -588173
rect 50 -587197 108 -587185
rect 50 -588173 62 -587197
rect 96 -588173 108 -587197
rect 50 -588185 108 -588173
rect -108 -588415 -50 -588403
rect -108 -589391 -96 -588415
rect -62 -589391 -50 -588415
rect -108 -589403 -50 -589391
rect 50 -588415 108 -588403
rect 50 -589391 62 -588415
rect 96 -589391 108 -588415
rect 50 -589403 108 -589391
rect -108 -589633 -50 -589621
rect -108 -590609 -96 -589633
rect -62 -590609 -50 -589633
rect -108 -590621 -50 -590609
rect 50 -589633 108 -589621
rect 50 -590609 62 -589633
rect 96 -590609 108 -589633
rect 50 -590621 108 -590609
rect -108 -590851 -50 -590839
rect -108 -591827 -96 -590851
rect -62 -591827 -50 -590851
rect -108 -591839 -50 -591827
rect 50 -590851 108 -590839
rect 50 -591827 62 -590851
rect 96 -591827 108 -590851
rect 50 -591839 108 -591827
rect -108 -592069 -50 -592057
rect -108 -593045 -96 -592069
rect -62 -593045 -50 -592069
rect -108 -593057 -50 -593045
rect 50 -592069 108 -592057
rect 50 -593045 62 -592069
rect 96 -593045 108 -592069
rect 50 -593057 108 -593045
rect -108 -593287 -50 -593275
rect -108 -594263 -96 -593287
rect -62 -594263 -50 -593287
rect -108 -594275 -50 -594263
rect 50 -593287 108 -593275
rect 50 -594263 62 -593287
rect 96 -594263 108 -593287
rect 50 -594275 108 -594263
rect -108 -594505 -50 -594493
rect -108 -595481 -96 -594505
rect -62 -595481 -50 -594505
rect -108 -595493 -50 -595481
rect 50 -594505 108 -594493
rect 50 -595481 62 -594505
rect 96 -595481 108 -594505
rect 50 -595493 108 -595481
rect -108 -595723 -50 -595711
rect -108 -596699 -96 -595723
rect -62 -596699 -50 -595723
rect -108 -596711 -50 -596699
rect 50 -595723 108 -595711
rect 50 -596699 62 -595723
rect 96 -596699 108 -595723
rect 50 -596711 108 -596699
rect -108 -596941 -50 -596929
rect -108 -597917 -96 -596941
rect -62 -597917 -50 -596941
rect -108 -597929 -50 -597917
rect 50 -596941 108 -596929
rect 50 -597917 62 -596941
rect 96 -597917 108 -596941
rect 50 -597929 108 -597917
rect -108 -598159 -50 -598147
rect -108 -599135 -96 -598159
rect -62 -599135 -50 -598159
rect -108 -599147 -50 -599135
rect 50 -598159 108 -598147
rect 50 -599135 62 -598159
rect 96 -599135 108 -598159
rect 50 -599147 108 -599135
rect -108 -599377 -50 -599365
rect -108 -600353 -96 -599377
rect -62 -600353 -50 -599377
rect -108 -600365 -50 -600353
rect 50 -599377 108 -599365
rect 50 -600353 62 -599377
rect 96 -600353 108 -599377
rect 50 -600365 108 -600353
rect -108 -600595 -50 -600583
rect -108 -601571 -96 -600595
rect -62 -601571 -50 -600595
rect -108 -601583 -50 -601571
rect 50 -600595 108 -600583
rect 50 -601571 62 -600595
rect 96 -601571 108 -600595
rect 50 -601583 108 -601571
rect -108 -601813 -50 -601801
rect -108 -602789 -96 -601813
rect -62 -602789 -50 -601813
rect -108 -602801 -50 -602789
rect 50 -601813 108 -601801
rect 50 -602789 62 -601813
rect 96 -602789 108 -601813
rect 50 -602801 108 -602789
rect -108 -603031 -50 -603019
rect -108 -604007 -96 -603031
rect -62 -604007 -50 -603031
rect -108 -604019 -50 -604007
rect 50 -603031 108 -603019
rect 50 -604007 62 -603031
rect 96 -604007 108 -603031
rect 50 -604019 108 -604007
rect -108 -604249 -50 -604237
rect -108 -605225 -96 -604249
rect -62 -605225 -50 -604249
rect -108 -605237 -50 -605225
rect 50 -604249 108 -604237
rect 50 -605225 62 -604249
rect 96 -605225 108 -604249
rect 50 -605237 108 -605225
rect -108 -605467 -50 -605455
rect -108 -606443 -96 -605467
rect -62 -606443 -50 -605467
rect -108 -606455 -50 -606443
rect 50 -605467 108 -605455
rect 50 -606443 62 -605467
rect 96 -606443 108 -605467
rect 50 -606455 108 -606443
rect -108 -606685 -50 -606673
rect -108 -607661 -96 -606685
rect -62 -607661 -50 -606685
rect -108 -607673 -50 -607661
rect 50 -606685 108 -606673
rect 50 -607661 62 -606685
rect 96 -607661 108 -606685
rect 50 -607673 108 -607661
rect -108 -607903 -50 -607891
rect -108 -608879 -96 -607903
rect -62 -608879 -50 -607903
rect -108 -608891 -50 -608879
rect 50 -607903 108 -607891
rect 50 -608879 62 -607903
rect 96 -608879 108 -607903
rect 50 -608891 108 -608879
<< mvndiffc >>
rect -96 607903 -62 608879
rect 62 607903 96 608879
rect -96 606685 -62 607661
rect 62 606685 96 607661
rect -96 605467 -62 606443
rect 62 605467 96 606443
rect -96 604249 -62 605225
rect 62 604249 96 605225
rect -96 603031 -62 604007
rect 62 603031 96 604007
rect -96 601813 -62 602789
rect 62 601813 96 602789
rect -96 600595 -62 601571
rect 62 600595 96 601571
rect -96 599377 -62 600353
rect 62 599377 96 600353
rect -96 598159 -62 599135
rect 62 598159 96 599135
rect -96 596941 -62 597917
rect 62 596941 96 597917
rect -96 595723 -62 596699
rect 62 595723 96 596699
rect -96 594505 -62 595481
rect 62 594505 96 595481
rect -96 593287 -62 594263
rect 62 593287 96 594263
rect -96 592069 -62 593045
rect 62 592069 96 593045
rect -96 590851 -62 591827
rect 62 590851 96 591827
rect -96 589633 -62 590609
rect 62 589633 96 590609
rect -96 588415 -62 589391
rect 62 588415 96 589391
rect -96 587197 -62 588173
rect 62 587197 96 588173
rect -96 585979 -62 586955
rect 62 585979 96 586955
rect -96 584761 -62 585737
rect 62 584761 96 585737
rect -96 583543 -62 584519
rect 62 583543 96 584519
rect -96 582325 -62 583301
rect 62 582325 96 583301
rect -96 581107 -62 582083
rect 62 581107 96 582083
rect -96 579889 -62 580865
rect 62 579889 96 580865
rect -96 578671 -62 579647
rect 62 578671 96 579647
rect -96 577453 -62 578429
rect 62 577453 96 578429
rect -96 576235 -62 577211
rect 62 576235 96 577211
rect -96 575017 -62 575993
rect 62 575017 96 575993
rect -96 573799 -62 574775
rect 62 573799 96 574775
rect -96 572581 -62 573557
rect 62 572581 96 573557
rect -96 571363 -62 572339
rect 62 571363 96 572339
rect -96 570145 -62 571121
rect 62 570145 96 571121
rect -96 568927 -62 569903
rect 62 568927 96 569903
rect -96 567709 -62 568685
rect 62 567709 96 568685
rect -96 566491 -62 567467
rect 62 566491 96 567467
rect -96 565273 -62 566249
rect 62 565273 96 566249
rect -96 564055 -62 565031
rect 62 564055 96 565031
rect -96 562837 -62 563813
rect 62 562837 96 563813
rect -96 561619 -62 562595
rect 62 561619 96 562595
rect -96 560401 -62 561377
rect 62 560401 96 561377
rect -96 559183 -62 560159
rect 62 559183 96 560159
rect -96 557965 -62 558941
rect 62 557965 96 558941
rect -96 556747 -62 557723
rect 62 556747 96 557723
rect -96 555529 -62 556505
rect 62 555529 96 556505
rect -96 554311 -62 555287
rect 62 554311 96 555287
rect -96 553093 -62 554069
rect 62 553093 96 554069
rect -96 551875 -62 552851
rect 62 551875 96 552851
rect -96 550657 -62 551633
rect 62 550657 96 551633
rect -96 549439 -62 550415
rect 62 549439 96 550415
rect -96 548221 -62 549197
rect 62 548221 96 549197
rect -96 547003 -62 547979
rect 62 547003 96 547979
rect -96 545785 -62 546761
rect 62 545785 96 546761
rect -96 544567 -62 545543
rect 62 544567 96 545543
rect -96 543349 -62 544325
rect 62 543349 96 544325
rect -96 542131 -62 543107
rect 62 542131 96 543107
rect -96 540913 -62 541889
rect 62 540913 96 541889
rect -96 539695 -62 540671
rect 62 539695 96 540671
rect -96 538477 -62 539453
rect 62 538477 96 539453
rect -96 537259 -62 538235
rect 62 537259 96 538235
rect -96 536041 -62 537017
rect 62 536041 96 537017
rect -96 534823 -62 535799
rect 62 534823 96 535799
rect -96 533605 -62 534581
rect 62 533605 96 534581
rect -96 532387 -62 533363
rect 62 532387 96 533363
rect -96 531169 -62 532145
rect 62 531169 96 532145
rect -96 529951 -62 530927
rect 62 529951 96 530927
rect -96 528733 -62 529709
rect 62 528733 96 529709
rect -96 527515 -62 528491
rect 62 527515 96 528491
rect -96 526297 -62 527273
rect 62 526297 96 527273
rect -96 525079 -62 526055
rect 62 525079 96 526055
rect -96 523861 -62 524837
rect 62 523861 96 524837
rect -96 522643 -62 523619
rect 62 522643 96 523619
rect -96 521425 -62 522401
rect 62 521425 96 522401
rect -96 520207 -62 521183
rect 62 520207 96 521183
rect -96 518989 -62 519965
rect 62 518989 96 519965
rect -96 517771 -62 518747
rect 62 517771 96 518747
rect -96 516553 -62 517529
rect 62 516553 96 517529
rect -96 515335 -62 516311
rect 62 515335 96 516311
rect -96 514117 -62 515093
rect 62 514117 96 515093
rect -96 512899 -62 513875
rect 62 512899 96 513875
rect -96 511681 -62 512657
rect 62 511681 96 512657
rect -96 510463 -62 511439
rect 62 510463 96 511439
rect -96 509245 -62 510221
rect 62 509245 96 510221
rect -96 508027 -62 509003
rect 62 508027 96 509003
rect -96 506809 -62 507785
rect 62 506809 96 507785
rect -96 505591 -62 506567
rect 62 505591 96 506567
rect -96 504373 -62 505349
rect 62 504373 96 505349
rect -96 503155 -62 504131
rect 62 503155 96 504131
rect -96 501937 -62 502913
rect 62 501937 96 502913
rect -96 500719 -62 501695
rect 62 500719 96 501695
rect -96 499501 -62 500477
rect 62 499501 96 500477
rect -96 498283 -62 499259
rect 62 498283 96 499259
rect -96 497065 -62 498041
rect 62 497065 96 498041
rect -96 495847 -62 496823
rect 62 495847 96 496823
rect -96 494629 -62 495605
rect 62 494629 96 495605
rect -96 493411 -62 494387
rect 62 493411 96 494387
rect -96 492193 -62 493169
rect 62 492193 96 493169
rect -96 490975 -62 491951
rect 62 490975 96 491951
rect -96 489757 -62 490733
rect 62 489757 96 490733
rect -96 488539 -62 489515
rect 62 488539 96 489515
rect -96 487321 -62 488297
rect 62 487321 96 488297
rect -96 486103 -62 487079
rect 62 486103 96 487079
rect -96 484885 -62 485861
rect 62 484885 96 485861
rect -96 483667 -62 484643
rect 62 483667 96 484643
rect -96 482449 -62 483425
rect 62 482449 96 483425
rect -96 481231 -62 482207
rect 62 481231 96 482207
rect -96 480013 -62 480989
rect 62 480013 96 480989
rect -96 478795 -62 479771
rect 62 478795 96 479771
rect -96 477577 -62 478553
rect 62 477577 96 478553
rect -96 476359 -62 477335
rect 62 476359 96 477335
rect -96 475141 -62 476117
rect 62 475141 96 476117
rect -96 473923 -62 474899
rect 62 473923 96 474899
rect -96 472705 -62 473681
rect 62 472705 96 473681
rect -96 471487 -62 472463
rect 62 471487 96 472463
rect -96 470269 -62 471245
rect 62 470269 96 471245
rect -96 469051 -62 470027
rect 62 469051 96 470027
rect -96 467833 -62 468809
rect 62 467833 96 468809
rect -96 466615 -62 467591
rect 62 466615 96 467591
rect -96 465397 -62 466373
rect 62 465397 96 466373
rect -96 464179 -62 465155
rect 62 464179 96 465155
rect -96 462961 -62 463937
rect 62 462961 96 463937
rect -96 461743 -62 462719
rect 62 461743 96 462719
rect -96 460525 -62 461501
rect 62 460525 96 461501
rect -96 459307 -62 460283
rect 62 459307 96 460283
rect -96 458089 -62 459065
rect 62 458089 96 459065
rect -96 456871 -62 457847
rect 62 456871 96 457847
rect -96 455653 -62 456629
rect 62 455653 96 456629
rect -96 454435 -62 455411
rect 62 454435 96 455411
rect -96 453217 -62 454193
rect 62 453217 96 454193
rect -96 451999 -62 452975
rect 62 451999 96 452975
rect -96 450781 -62 451757
rect 62 450781 96 451757
rect -96 449563 -62 450539
rect 62 449563 96 450539
rect -96 448345 -62 449321
rect 62 448345 96 449321
rect -96 447127 -62 448103
rect 62 447127 96 448103
rect -96 445909 -62 446885
rect 62 445909 96 446885
rect -96 444691 -62 445667
rect 62 444691 96 445667
rect -96 443473 -62 444449
rect 62 443473 96 444449
rect -96 442255 -62 443231
rect 62 442255 96 443231
rect -96 441037 -62 442013
rect 62 441037 96 442013
rect -96 439819 -62 440795
rect 62 439819 96 440795
rect -96 438601 -62 439577
rect 62 438601 96 439577
rect -96 437383 -62 438359
rect 62 437383 96 438359
rect -96 436165 -62 437141
rect 62 436165 96 437141
rect -96 434947 -62 435923
rect 62 434947 96 435923
rect -96 433729 -62 434705
rect 62 433729 96 434705
rect -96 432511 -62 433487
rect 62 432511 96 433487
rect -96 431293 -62 432269
rect 62 431293 96 432269
rect -96 430075 -62 431051
rect 62 430075 96 431051
rect -96 428857 -62 429833
rect 62 428857 96 429833
rect -96 427639 -62 428615
rect 62 427639 96 428615
rect -96 426421 -62 427397
rect 62 426421 96 427397
rect -96 425203 -62 426179
rect 62 425203 96 426179
rect -96 423985 -62 424961
rect 62 423985 96 424961
rect -96 422767 -62 423743
rect 62 422767 96 423743
rect -96 421549 -62 422525
rect 62 421549 96 422525
rect -96 420331 -62 421307
rect 62 420331 96 421307
rect -96 419113 -62 420089
rect 62 419113 96 420089
rect -96 417895 -62 418871
rect 62 417895 96 418871
rect -96 416677 -62 417653
rect 62 416677 96 417653
rect -96 415459 -62 416435
rect 62 415459 96 416435
rect -96 414241 -62 415217
rect 62 414241 96 415217
rect -96 413023 -62 413999
rect 62 413023 96 413999
rect -96 411805 -62 412781
rect 62 411805 96 412781
rect -96 410587 -62 411563
rect 62 410587 96 411563
rect -96 409369 -62 410345
rect 62 409369 96 410345
rect -96 408151 -62 409127
rect 62 408151 96 409127
rect -96 406933 -62 407909
rect 62 406933 96 407909
rect -96 405715 -62 406691
rect 62 405715 96 406691
rect -96 404497 -62 405473
rect 62 404497 96 405473
rect -96 403279 -62 404255
rect 62 403279 96 404255
rect -96 402061 -62 403037
rect 62 402061 96 403037
rect -96 400843 -62 401819
rect 62 400843 96 401819
rect -96 399625 -62 400601
rect 62 399625 96 400601
rect -96 398407 -62 399383
rect 62 398407 96 399383
rect -96 397189 -62 398165
rect 62 397189 96 398165
rect -96 395971 -62 396947
rect 62 395971 96 396947
rect -96 394753 -62 395729
rect 62 394753 96 395729
rect -96 393535 -62 394511
rect 62 393535 96 394511
rect -96 392317 -62 393293
rect 62 392317 96 393293
rect -96 391099 -62 392075
rect 62 391099 96 392075
rect -96 389881 -62 390857
rect 62 389881 96 390857
rect -96 388663 -62 389639
rect 62 388663 96 389639
rect -96 387445 -62 388421
rect 62 387445 96 388421
rect -96 386227 -62 387203
rect 62 386227 96 387203
rect -96 385009 -62 385985
rect 62 385009 96 385985
rect -96 383791 -62 384767
rect 62 383791 96 384767
rect -96 382573 -62 383549
rect 62 382573 96 383549
rect -96 381355 -62 382331
rect 62 381355 96 382331
rect -96 380137 -62 381113
rect 62 380137 96 381113
rect -96 378919 -62 379895
rect 62 378919 96 379895
rect -96 377701 -62 378677
rect 62 377701 96 378677
rect -96 376483 -62 377459
rect 62 376483 96 377459
rect -96 375265 -62 376241
rect 62 375265 96 376241
rect -96 374047 -62 375023
rect 62 374047 96 375023
rect -96 372829 -62 373805
rect 62 372829 96 373805
rect -96 371611 -62 372587
rect 62 371611 96 372587
rect -96 370393 -62 371369
rect 62 370393 96 371369
rect -96 369175 -62 370151
rect 62 369175 96 370151
rect -96 367957 -62 368933
rect 62 367957 96 368933
rect -96 366739 -62 367715
rect 62 366739 96 367715
rect -96 365521 -62 366497
rect 62 365521 96 366497
rect -96 364303 -62 365279
rect 62 364303 96 365279
rect -96 363085 -62 364061
rect 62 363085 96 364061
rect -96 361867 -62 362843
rect 62 361867 96 362843
rect -96 360649 -62 361625
rect 62 360649 96 361625
rect -96 359431 -62 360407
rect 62 359431 96 360407
rect -96 358213 -62 359189
rect 62 358213 96 359189
rect -96 356995 -62 357971
rect 62 356995 96 357971
rect -96 355777 -62 356753
rect 62 355777 96 356753
rect -96 354559 -62 355535
rect 62 354559 96 355535
rect -96 353341 -62 354317
rect 62 353341 96 354317
rect -96 352123 -62 353099
rect 62 352123 96 353099
rect -96 350905 -62 351881
rect 62 350905 96 351881
rect -96 349687 -62 350663
rect 62 349687 96 350663
rect -96 348469 -62 349445
rect 62 348469 96 349445
rect -96 347251 -62 348227
rect 62 347251 96 348227
rect -96 346033 -62 347009
rect 62 346033 96 347009
rect -96 344815 -62 345791
rect 62 344815 96 345791
rect -96 343597 -62 344573
rect 62 343597 96 344573
rect -96 342379 -62 343355
rect 62 342379 96 343355
rect -96 341161 -62 342137
rect 62 341161 96 342137
rect -96 339943 -62 340919
rect 62 339943 96 340919
rect -96 338725 -62 339701
rect 62 338725 96 339701
rect -96 337507 -62 338483
rect 62 337507 96 338483
rect -96 336289 -62 337265
rect 62 336289 96 337265
rect -96 335071 -62 336047
rect 62 335071 96 336047
rect -96 333853 -62 334829
rect 62 333853 96 334829
rect -96 332635 -62 333611
rect 62 332635 96 333611
rect -96 331417 -62 332393
rect 62 331417 96 332393
rect -96 330199 -62 331175
rect 62 330199 96 331175
rect -96 328981 -62 329957
rect 62 328981 96 329957
rect -96 327763 -62 328739
rect 62 327763 96 328739
rect -96 326545 -62 327521
rect 62 326545 96 327521
rect -96 325327 -62 326303
rect 62 325327 96 326303
rect -96 324109 -62 325085
rect 62 324109 96 325085
rect -96 322891 -62 323867
rect 62 322891 96 323867
rect -96 321673 -62 322649
rect 62 321673 96 322649
rect -96 320455 -62 321431
rect 62 320455 96 321431
rect -96 319237 -62 320213
rect 62 319237 96 320213
rect -96 318019 -62 318995
rect 62 318019 96 318995
rect -96 316801 -62 317777
rect 62 316801 96 317777
rect -96 315583 -62 316559
rect 62 315583 96 316559
rect -96 314365 -62 315341
rect 62 314365 96 315341
rect -96 313147 -62 314123
rect 62 313147 96 314123
rect -96 311929 -62 312905
rect 62 311929 96 312905
rect -96 310711 -62 311687
rect 62 310711 96 311687
rect -96 309493 -62 310469
rect 62 309493 96 310469
rect -96 308275 -62 309251
rect 62 308275 96 309251
rect -96 307057 -62 308033
rect 62 307057 96 308033
rect -96 305839 -62 306815
rect 62 305839 96 306815
rect -96 304621 -62 305597
rect 62 304621 96 305597
rect -96 303403 -62 304379
rect 62 303403 96 304379
rect -96 302185 -62 303161
rect 62 302185 96 303161
rect -96 300967 -62 301943
rect 62 300967 96 301943
rect -96 299749 -62 300725
rect 62 299749 96 300725
rect -96 298531 -62 299507
rect 62 298531 96 299507
rect -96 297313 -62 298289
rect 62 297313 96 298289
rect -96 296095 -62 297071
rect 62 296095 96 297071
rect -96 294877 -62 295853
rect 62 294877 96 295853
rect -96 293659 -62 294635
rect 62 293659 96 294635
rect -96 292441 -62 293417
rect 62 292441 96 293417
rect -96 291223 -62 292199
rect 62 291223 96 292199
rect -96 290005 -62 290981
rect 62 290005 96 290981
rect -96 288787 -62 289763
rect 62 288787 96 289763
rect -96 287569 -62 288545
rect 62 287569 96 288545
rect -96 286351 -62 287327
rect 62 286351 96 287327
rect -96 285133 -62 286109
rect 62 285133 96 286109
rect -96 283915 -62 284891
rect 62 283915 96 284891
rect -96 282697 -62 283673
rect 62 282697 96 283673
rect -96 281479 -62 282455
rect 62 281479 96 282455
rect -96 280261 -62 281237
rect 62 280261 96 281237
rect -96 279043 -62 280019
rect 62 279043 96 280019
rect -96 277825 -62 278801
rect 62 277825 96 278801
rect -96 276607 -62 277583
rect 62 276607 96 277583
rect -96 275389 -62 276365
rect 62 275389 96 276365
rect -96 274171 -62 275147
rect 62 274171 96 275147
rect -96 272953 -62 273929
rect 62 272953 96 273929
rect -96 271735 -62 272711
rect 62 271735 96 272711
rect -96 270517 -62 271493
rect 62 270517 96 271493
rect -96 269299 -62 270275
rect 62 269299 96 270275
rect -96 268081 -62 269057
rect 62 268081 96 269057
rect -96 266863 -62 267839
rect 62 266863 96 267839
rect -96 265645 -62 266621
rect 62 265645 96 266621
rect -96 264427 -62 265403
rect 62 264427 96 265403
rect -96 263209 -62 264185
rect 62 263209 96 264185
rect -96 261991 -62 262967
rect 62 261991 96 262967
rect -96 260773 -62 261749
rect 62 260773 96 261749
rect -96 259555 -62 260531
rect 62 259555 96 260531
rect -96 258337 -62 259313
rect 62 258337 96 259313
rect -96 257119 -62 258095
rect 62 257119 96 258095
rect -96 255901 -62 256877
rect 62 255901 96 256877
rect -96 254683 -62 255659
rect 62 254683 96 255659
rect -96 253465 -62 254441
rect 62 253465 96 254441
rect -96 252247 -62 253223
rect 62 252247 96 253223
rect -96 251029 -62 252005
rect 62 251029 96 252005
rect -96 249811 -62 250787
rect 62 249811 96 250787
rect -96 248593 -62 249569
rect 62 248593 96 249569
rect -96 247375 -62 248351
rect 62 247375 96 248351
rect -96 246157 -62 247133
rect 62 246157 96 247133
rect -96 244939 -62 245915
rect 62 244939 96 245915
rect -96 243721 -62 244697
rect 62 243721 96 244697
rect -96 242503 -62 243479
rect 62 242503 96 243479
rect -96 241285 -62 242261
rect 62 241285 96 242261
rect -96 240067 -62 241043
rect 62 240067 96 241043
rect -96 238849 -62 239825
rect 62 238849 96 239825
rect -96 237631 -62 238607
rect 62 237631 96 238607
rect -96 236413 -62 237389
rect 62 236413 96 237389
rect -96 235195 -62 236171
rect 62 235195 96 236171
rect -96 233977 -62 234953
rect 62 233977 96 234953
rect -96 232759 -62 233735
rect 62 232759 96 233735
rect -96 231541 -62 232517
rect 62 231541 96 232517
rect -96 230323 -62 231299
rect 62 230323 96 231299
rect -96 229105 -62 230081
rect 62 229105 96 230081
rect -96 227887 -62 228863
rect 62 227887 96 228863
rect -96 226669 -62 227645
rect 62 226669 96 227645
rect -96 225451 -62 226427
rect 62 225451 96 226427
rect -96 224233 -62 225209
rect 62 224233 96 225209
rect -96 223015 -62 223991
rect 62 223015 96 223991
rect -96 221797 -62 222773
rect 62 221797 96 222773
rect -96 220579 -62 221555
rect 62 220579 96 221555
rect -96 219361 -62 220337
rect 62 219361 96 220337
rect -96 218143 -62 219119
rect 62 218143 96 219119
rect -96 216925 -62 217901
rect 62 216925 96 217901
rect -96 215707 -62 216683
rect 62 215707 96 216683
rect -96 214489 -62 215465
rect 62 214489 96 215465
rect -96 213271 -62 214247
rect 62 213271 96 214247
rect -96 212053 -62 213029
rect 62 212053 96 213029
rect -96 210835 -62 211811
rect 62 210835 96 211811
rect -96 209617 -62 210593
rect 62 209617 96 210593
rect -96 208399 -62 209375
rect 62 208399 96 209375
rect -96 207181 -62 208157
rect 62 207181 96 208157
rect -96 205963 -62 206939
rect 62 205963 96 206939
rect -96 204745 -62 205721
rect 62 204745 96 205721
rect -96 203527 -62 204503
rect 62 203527 96 204503
rect -96 202309 -62 203285
rect 62 202309 96 203285
rect -96 201091 -62 202067
rect 62 201091 96 202067
rect -96 199873 -62 200849
rect 62 199873 96 200849
rect -96 198655 -62 199631
rect 62 198655 96 199631
rect -96 197437 -62 198413
rect 62 197437 96 198413
rect -96 196219 -62 197195
rect 62 196219 96 197195
rect -96 195001 -62 195977
rect 62 195001 96 195977
rect -96 193783 -62 194759
rect 62 193783 96 194759
rect -96 192565 -62 193541
rect 62 192565 96 193541
rect -96 191347 -62 192323
rect 62 191347 96 192323
rect -96 190129 -62 191105
rect 62 190129 96 191105
rect -96 188911 -62 189887
rect 62 188911 96 189887
rect -96 187693 -62 188669
rect 62 187693 96 188669
rect -96 186475 -62 187451
rect 62 186475 96 187451
rect -96 185257 -62 186233
rect 62 185257 96 186233
rect -96 184039 -62 185015
rect 62 184039 96 185015
rect -96 182821 -62 183797
rect 62 182821 96 183797
rect -96 181603 -62 182579
rect 62 181603 96 182579
rect -96 180385 -62 181361
rect 62 180385 96 181361
rect -96 179167 -62 180143
rect 62 179167 96 180143
rect -96 177949 -62 178925
rect 62 177949 96 178925
rect -96 176731 -62 177707
rect 62 176731 96 177707
rect -96 175513 -62 176489
rect 62 175513 96 176489
rect -96 174295 -62 175271
rect 62 174295 96 175271
rect -96 173077 -62 174053
rect 62 173077 96 174053
rect -96 171859 -62 172835
rect 62 171859 96 172835
rect -96 170641 -62 171617
rect 62 170641 96 171617
rect -96 169423 -62 170399
rect 62 169423 96 170399
rect -96 168205 -62 169181
rect 62 168205 96 169181
rect -96 166987 -62 167963
rect 62 166987 96 167963
rect -96 165769 -62 166745
rect 62 165769 96 166745
rect -96 164551 -62 165527
rect 62 164551 96 165527
rect -96 163333 -62 164309
rect 62 163333 96 164309
rect -96 162115 -62 163091
rect 62 162115 96 163091
rect -96 160897 -62 161873
rect 62 160897 96 161873
rect -96 159679 -62 160655
rect 62 159679 96 160655
rect -96 158461 -62 159437
rect 62 158461 96 159437
rect -96 157243 -62 158219
rect 62 157243 96 158219
rect -96 156025 -62 157001
rect 62 156025 96 157001
rect -96 154807 -62 155783
rect 62 154807 96 155783
rect -96 153589 -62 154565
rect 62 153589 96 154565
rect -96 152371 -62 153347
rect 62 152371 96 153347
rect -96 151153 -62 152129
rect 62 151153 96 152129
rect -96 149935 -62 150911
rect 62 149935 96 150911
rect -96 148717 -62 149693
rect 62 148717 96 149693
rect -96 147499 -62 148475
rect 62 147499 96 148475
rect -96 146281 -62 147257
rect 62 146281 96 147257
rect -96 145063 -62 146039
rect 62 145063 96 146039
rect -96 143845 -62 144821
rect 62 143845 96 144821
rect -96 142627 -62 143603
rect 62 142627 96 143603
rect -96 141409 -62 142385
rect 62 141409 96 142385
rect -96 140191 -62 141167
rect 62 140191 96 141167
rect -96 138973 -62 139949
rect 62 138973 96 139949
rect -96 137755 -62 138731
rect 62 137755 96 138731
rect -96 136537 -62 137513
rect 62 136537 96 137513
rect -96 135319 -62 136295
rect 62 135319 96 136295
rect -96 134101 -62 135077
rect 62 134101 96 135077
rect -96 132883 -62 133859
rect 62 132883 96 133859
rect -96 131665 -62 132641
rect 62 131665 96 132641
rect -96 130447 -62 131423
rect 62 130447 96 131423
rect -96 129229 -62 130205
rect 62 129229 96 130205
rect -96 128011 -62 128987
rect 62 128011 96 128987
rect -96 126793 -62 127769
rect 62 126793 96 127769
rect -96 125575 -62 126551
rect 62 125575 96 126551
rect -96 124357 -62 125333
rect 62 124357 96 125333
rect -96 123139 -62 124115
rect 62 123139 96 124115
rect -96 121921 -62 122897
rect 62 121921 96 122897
rect -96 120703 -62 121679
rect 62 120703 96 121679
rect -96 119485 -62 120461
rect 62 119485 96 120461
rect -96 118267 -62 119243
rect 62 118267 96 119243
rect -96 117049 -62 118025
rect 62 117049 96 118025
rect -96 115831 -62 116807
rect 62 115831 96 116807
rect -96 114613 -62 115589
rect 62 114613 96 115589
rect -96 113395 -62 114371
rect 62 113395 96 114371
rect -96 112177 -62 113153
rect 62 112177 96 113153
rect -96 110959 -62 111935
rect 62 110959 96 111935
rect -96 109741 -62 110717
rect 62 109741 96 110717
rect -96 108523 -62 109499
rect 62 108523 96 109499
rect -96 107305 -62 108281
rect 62 107305 96 108281
rect -96 106087 -62 107063
rect 62 106087 96 107063
rect -96 104869 -62 105845
rect 62 104869 96 105845
rect -96 103651 -62 104627
rect 62 103651 96 104627
rect -96 102433 -62 103409
rect 62 102433 96 103409
rect -96 101215 -62 102191
rect 62 101215 96 102191
rect -96 99997 -62 100973
rect 62 99997 96 100973
rect -96 98779 -62 99755
rect 62 98779 96 99755
rect -96 97561 -62 98537
rect 62 97561 96 98537
rect -96 96343 -62 97319
rect 62 96343 96 97319
rect -96 95125 -62 96101
rect 62 95125 96 96101
rect -96 93907 -62 94883
rect 62 93907 96 94883
rect -96 92689 -62 93665
rect 62 92689 96 93665
rect -96 91471 -62 92447
rect 62 91471 96 92447
rect -96 90253 -62 91229
rect 62 90253 96 91229
rect -96 89035 -62 90011
rect 62 89035 96 90011
rect -96 87817 -62 88793
rect 62 87817 96 88793
rect -96 86599 -62 87575
rect 62 86599 96 87575
rect -96 85381 -62 86357
rect 62 85381 96 86357
rect -96 84163 -62 85139
rect 62 84163 96 85139
rect -96 82945 -62 83921
rect 62 82945 96 83921
rect -96 81727 -62 82703
rect 62 81727 96 82703
rect -96 80509 -62 81485
rect 62 80509 96 81485
rect -96 79291 -62 80267
rect 62 79291 96 80267
rect -96 78073 -62 79049
rect 62 78073 96 79049
rect -96 76855 -62 77831
rect 62 76855 96 77831
rect -96 75637 -62 76613
rect 62 75637 96 76613
rect -96 74419 -62 75395
rect 62 74419 96 75395
rect -96 73201 -62 74177
rect 62 73201 96 74177
rect -96 71983 -62 72959
rect 62 71983 96 72959
rect -96 70765 -62 71741
rect 62 70765 96 71741
rect -96 69547 -62 70523
rect 62 69547 96 70523
rect -96 68329 -62 69305
rect 62 68329 96 69305
rect -96 67111 -62 68087
rect 62 67111 96 68087
rect -96 65893 -62 66869
rect 62 65893 96 66869
rect -96 64675 -62 65651
rect 62 64675 96 65651
rect -96 63457 -62 64433
rect 62 63457 96 64433
rect -96 62239 -62 63215
rect 62 62239 96 63215
rect -96 61021 -62 61997
rect 62 61021 96 61997
rect -96 59803 -62 60779
rect 62 59803 96 60779
rect -96 58585 -62 59561
rect 62 58585 96 59561
rect -96 57367 -62 58343
rect 62 57367 96 58343
rect -96 56149 -62 57125
rect 62 56149 96 57125
rect -96 54931 -62 55907
rect 62 54931 96 55907
rect -96 53713 -62 54689
rect 62 53713 96 54689
rect -96 52495 -62 53471
rect 62 52495 96 53471
rect -96 51277 -62 52253
rect 62 51277 96 52253
rect -96 50059 -62 51035
rect 62 50059 96 51035
rect -96 48841 -62 49817
rect 62 48841 96 49817
rect -96 47623 -62 48599
rect 62 47623 96 48599
rect -96 46405 -62 47381
rect 62 46405 96 47381
rect -96 45187 -62 46163
rect 62 45187 96 46163
rect -96 43969 -62 44945
rect 62 43969 96 44945
rect -96 42751 -62 43727
rect 62 42751 96 43727
rect -96 41533 -62 42509
rect 62 41533 96 42509
rect -96 40315 -62 41291
rect 62 40315 96 41291
rect -96 39097 -62 40073
rect 62 39097 96 40073
rect -96 37879 -62 38855
rect 62 37879 96 38855
rect -96 36661 -62 37637
rect 62 36661 96 37637
rect -96 35443 -62 36419
rect 62 35443 96 36419
rect -96 34225 -62 35201
rect 62 34225 96 35201
rect -96 33007 -62 33983
rect 62 33007 96 33983
rect -96 31789 -62 32765
rect 62 31789 96 32765
rect -96 30571 -62 31547
rect 62 30571 96 31547
rect -96 29353 -62 30329
rect 62 29353 96 30329
rect -96 28135 -62 29111
rect 62 28135 96 29111
rect -96 26917 -62 27893
rect 62 26917 96 27893
rect -96 25699 -62 26675
rect 62 25699 96 26675
rect -96 24481 -62 25457
rect 62 24481 96 25457
rect -96 23263 -62 24239
rect 62 23263 96 24239
rect -96 22045 -62 23021
rect 62 22045 96 23021
rect -96 20827 -62 21803
rect 62 20827 96 21803
rect -96 19609 -62 20585
rect 62 19609 96 20585
rect -96 18391 -62 19367
rect 62 18391 96 19367
rect -96 17173 -62 18149
rect 62 17173 96 18149
rect -96 15955 -62 16931
rect 62 15955 96 16931
rect -96 14737 -62 15713
rect 62 14737 96 15713
rect -96 13519 -62 14495
rect 62 13519 96 14495
rect -96 12301 -62 13277
rect 62 12301 96 13277
rect -96 11083 -62 12059
rect 62 11083 96 12059
rect -96 9865 -62 10841
rect 62 9865 96 10841
rect -96 8647 -62 9623
rect 62 8647 96 9623
rect -96 7429 -62 8405
rect 62 7429 96 8405
rect -96 6211 -62 7187
rect 62 6211 96 7187
rect -96 4993 -62 5969
rect 62 4993 96 5969
rect -96 3775 -62 4751
rect 62 3775 96 4751
rect -96 2557 -62 3533
rect 62 2557 96 3533
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -96 121 -62 1097
rect 62 121 96 1097
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
rect -96 -3533 -62 -2557
rect 62 -3533 96 -2557
rect -96 -4751 -62 -3775
rect 62 -4751 96 -3775
rect -96 -5969 -62 -4993
rect 62 -5969 96 -4993
rect -96 -7187 -62 -6211
rect 62 -7187 96 -6211
rect -96 -8405 -62 -7429
rect 62 -8405 96 -7429
rect -96 -9623 -62 -8647
rect 62 -9623 96 -8647
rect -96 -10841 -62 -9865
rect 62 -10841 96 -9865
rect -96 -12059 -62 -11083
rect 62 -12059 96 -11083
rect -96 -13277 -62 -12301
rect 62 -13277 96 -12301
rect -96 -14495 -62 -13519
rect 62 -14495 96 -13519
rect -96 -15713 -62 -14737
rect 62 -15713 96 -14737
rect -96 -16931 -62 -15955
rect 62 -16931 96 -15955
rect -96 -18149 -62 -17173
rect 62 -18149 96 -17173
rect -96 -19367 -62 -18391
rect 62 -19367 96 -18391
rect -96 -20585 -62 -19609
rect 62 -20585 96 -19609
rect -96 -21803 -62 -20827
rect 62 -21803 96 -20827
rect -96 -23021 -62 -22045
rect 62 -23021 96 -22045
rect -96 -24239 -62 -23263
rect 62 -24239 96 -23263
rect -96 -25457 -62 -24481
rect 62 -25457 96 -24481
rect -96 -26675 -62 -25699
rect 62 -26675 96 -25699
rect -96 -27893 -62 -26917
rect 62 -27893 96 -26917
rect -96 -29111 -62 -28135
rect 62 -29111 96 -28135
rect -96 -30329 -62 -29353
rect 62 -30329 96 -29353
rect -96 -31547 -62 -30571
rect 62 -31547 96 -30571
rect -96 -32765 -62 -31789
rect 62 -32765 96 -31789
rect -96 -33983 -62 -33007
rect 62 -33983 96 -33007
rect -96 -35201 -62 -34225
rect 62 -35201 96 -34225
rect -96 -36419 -62 -35443
rect 62 -36419 96 -35443
rect -96 -37637 -62 -36661
rect 62 -37637 96 -36661
rect -96 -38855 -62 -37879
rect 62 -38855 96 -37879
rect -96 -40073 -62 -39097
rect 62 -40073 96 -39097
rect -96 -41291 -62 -40315
rect 62 -41291 96 -40315
rect -96 -42509 -62 -41533
rect 62 -42509 96 -41533
rect -96 -43727 -62 -42751
rect 62 -43727 96 -42751
rect -96 -44945 -62 -43969
rect 62 -44945 96 -43969
rect -96 -46163 -62 -45187
rect 62 -46163 96 -45187
rect -96 -47381 -62 -46405
rect 62 -47381 96 -46405
rect -96 -48599 -62 -47623
rect 62 -48599 96 -47623
rect -96 -49817 -62 -48841
rect 62 -49817 96 -48841
rect -96 -51035 -62 -50059
rect 62 -51035 96 -50059
rect -96 -52253 -62 -51277
rect 62 -52253 96 -51277
rect -96 -53471 -62 -52495
rect 62 -53471 96 -52495
rect -96 -54689 -62 -53713
rect 62 -54689 96 -53713
rect -96 -55907 -62 -54931
rect 62 -55907 96 -54931
rect -96 -57125 -62 -56149
rect 62 -57125 96 -56149
rect -96 -58343 -62 -57367
rect 62 -58343 96 -57367
rect -96 -59561 -62 -58585
rect 62 -59561 96 -58585
rect -96 -60779 -62 -59803
rect 62 -60779 96 -59803
rect -96 -61997 -62 -61021
rect 62 -61997 96 -61021
rect -96 -63215 -62 -62239
rect 62 -63215 96 -62239
rect -96 -64433 -62 -63457
rect 62 -64433 96 -63457
rect -96 -65651 -62 -64675
rect 62 -65651 96 -64675
rect -96 -66869 -62 -65893
rect 62 -66869 96 -65893
rect -96 -68087 -62 -67111
rect 62 -68087 96 -67111
rect -96 -69305 -62 -68329
rect 62 -69305 96 -68329
rect -96 -70523 -62 -69547
rect 62 -70523 96 -69547
rect -96 -71741 -62 -70765
rect 62 -71741 96 -70765
rect -96 -72959 -62 -71983
rect 62 -72959 96 -71983
rect -96 -74177 -62 -73201
rect 62 -74177 96 -73201
rect -96 -75395 -62 -74419
rect 62 -75395 96 -74419
rect -96 -76613 -62 -75637
rect 62 -76613 96 -75637
rect -96 -77831 -62 -76855
rect 62 -77831 96 -76855
rect -96 -79049 -62 -78073
rect 62 -79049 96 -78073
rect -96 -80267 -62 -79291
rect 62 -80267 96 -79291
rect -96 -81485 -62 -80509
rect 62 -81485 96 -80509
rect -96 -82703 -62 -81727
rect 62 -82703 96 -81727
rect -96 -83921 -62 -82945
rect 62 -83921 96 -82945
rect -96 -85139 -62 -84163
rect 62 -85139 96 -84163
rect -96 -86357 -62 -85381
rect 62 -86357 96 -85381
rect -96 -87575 -62 -86599
rect 62 -87575 96 -86599
rect -96 -88793 -62 -87817
rect 62 -88793 96 -87817
rect -96 -90011 -62 -89035
rect 62 -90011 96 -89035
rect -96 -91229 -62 -90253
rect 62 -91229 96 -90253
rect -96 -92447 -62 -91471
rect 62 -92447 96 -91471
rect -96 -93665 -62 -92689
rect 62 -93665 96 -92689
rect -96 -94883 -62 -93907
rect 62 -94883 96 -93907
rect -96 -96101 -62 -95125
rect 62 -96101 96 -95125
rect -96 -97319 -62 -96343
rect 62 -97319 96 -96343
rect -96 -98537 -62 -97561
rect 62 -98537 96 -97561
rect -96 -99755 -62 -98779
rect 62 -99755 96 -98779
rect -96 -100973 -62 -99997
rect 62 -100973 96 -99997
rect -96 -102191 -62 -101215
rect 62 -102191 96 -101215
rect -96 -103409 -62 -102433
rect 62 -103409 96 -102433
rect -96 -104627 -62 -103651
rect 62 -104627 96 -103651
rect -96 -105845 -62 -104869
rect 62 -105845 96 -104869
rect -96 -107063 -62 -106087
rect 62 -107063 96 -106087
rect -96 -108281 -62 -107305
rect 62 -108281 96 -107305
rect -96 -109499 -62 -108523
rect 62 -109499 96 -108523
rect -96 -110717 -62 -109741
rect 62 -110717 96 -109741
rect -96 -111935 -62 -110959
rect 62 -111935 96 -110959
rect -96 -113153 -62 -112177
rect 62 -113153 96 -112177
rect -96 -114371 -62 -113395
rect 62 -114371 96 -113395
rect -96 -115589 -62 -114613
rect 62 -115589 96 -114613
rect -96 -116807 -62 -115831
rect 62 -116807 96 -115831
rect -96 -118025 -62 -117049
rect 62 -118025 96 -117049
rect -96 -119243 -62 -118267
rect 62 -119243 96 -118267
rect -96 -120461 -62 -119485
rect 62 -120461 96 -119485
rect -96 -121679 -62 -120703
rect 62 -121679 96 -120703
rect -96 -122897 -62 -121921
rect 62 -122897 96 -121921
rect -96 -124115 -62 -123139
rect 62 -124115 96 -123139
rect -96 -125333 -62 -124357
rect 62 -125333 96 -124357
rect -96 -126551 -62 -125575
rect 62 -126551 96 -125575
rect -96 -127769 -62 -126793
rect 62 -127769 96 -126793
rect -96 -128987 -62 -128011
rect 62 -128987 96 -128011
rect -96 -130205 -62 -129229
rect 62 -130205 96 -129229
rect -96 -131423 -62 -130447
rect 62 -131423 96 -130447
rect -96 -132641 -62 -131665
rect 62 -132641 96 -131665
rect -96 -133859 -62 -132883
rect 62 -133859 96 -132883
rect -96 -135077 -62 -134101
rect 62 -135077 96 -134101
rect -96 -136295 -62 -135319
rect 62 -136295 96 -135319
rect -96 -137513 -62 -136537
rect 62 -137513 96 -136537
rect -96 -138731 -62 -137755
rect 62 -138731 96 -137755
rect -96 -139949 -62 -138973
rect 62 -139949 96 -138973
rect -96 -141167 -62 -140191
rect 62 -141167 96 -140191
rect -96 -142385 -62 -141409
rect 62 -142385 96 -141409
rect -96 -143603 -62 -142627
rect 62 -143603 96 -142627
rect -96 -144821 -62 -143845
rect 62 -144821 96 -143845
rect -96 -146039 -62 -145063
rect 62 -146039 96 -145063
rect -96 -147257 -62 -146281
rect 62 -147257 96 -146281
rect -96 -148475 -62 -147499
rect 62 -148475 96 -147499
rect -96 -149693 -62 -148717
rect 62 -149693 96 -148717
rect -96 -150911 -62 -149935
rect 62 -150911 96 -149935
rect -96 -152129 -62 -151153
rect 62 -152129 96 -151153
rect -96 -153347 -62 -152371
rect 62 -153347 96 -152371
rect -96 -154565 -62 -153589
rect 62 -154565 96 -153589
rect -96 -155783 -62 -154807
rect 62 -155783 96 -154807
rect -96 -157001 -62 -156025
rect 62 -157001 96 -156025
rect -96 -158219 -62 -157243
rect 62 -158219 96 -157243
rect -96 -159437 -62 -158461
rect 62 -159437 96 -158461
rect -96 -160655 -62 -159679
rect 62 -160655 96 -159679
rect -96 -161873 -62 -160897
rect 62 -161873 96 -160897
rect -96 -163091 -62 -162115
rect 62 -163091 96 -162115
rect -96 -164309 -62 -163333
rect 62 -164309 96 -163333
rect -96 -165527 -62 -164551
rect 62 -165527 96 -164551
rect -96 -166745 -62 -165769
rect 62 -166745 96 -165769
rect -96 -167963 -62 -166987
rect 62 -167963 96 -166987
rect -96 -169181 -62 -168205
rect 62 -169181 96 -168205
rect -96 -170399 -62 -169423
rect 62 -170399 96 -169423
rect -96 -171617 -62 -170641
rect 62 -171617 96 -170641
rect -96 -172835 -62 -171859
rect 62 -172835 96 -171859
rect -96 -174053 -62 -173077
rect 62 -174053 96 -173077
rect -96 -175271 -62 -174295
rect 62 -175271 96 -174295
rect -96 -176489 -62 -175513
rect 62 -176489 96 -175513
rect -96 -177707 -62 -176731
rect 62 -177707 96 -176731
rect -96 -178925 -62 -177949
rect 62 -178925 96 -177949
rect -96 -180143 -62 -179167
rect 62 -180143 96 -179167
rect -96 -181361 -62 -180385
rect 62 -181361 96 -180385
rect -96 -182579 -62 -181603
rect 62 -182579 96 -181603
rect -96 -183797 -62 -182821
rect 62 -183797 96 -182821
rect -96 -185015 -62 -184039
rect 62 -185015 96 -184039
rect -96 -186233 -62 -185257
rect 62 -186233 96 -185257
rect -96 -187451 -62 -186475
rect 62 -187451 96 -186475
rect -96 -188669 -62 -187693
rect 62 -188669 96 -187693
rect -96 -189887 -62 -188911
rect 62 -189887 96 -188911
rect -96 -191105 -62 -190129
rect 62 -191105 96 -190129
rect -96 -192323 -62 -191347
rect 62 -192323 96 -191347
rect -96 -193541 -62 -192565
rect 62 -193541 96 -192565
rect -96 -194759 -62 -193783
rect 62 -194759 96 -193783
rect -96 -195977 -62 -195001
rect 62 -195977 96 -195001
rect -96 -197195 -62 -196219
rect 62 -197195 96 -196219
rect -96 -198413 -62 -197437
rect 62 -198413 96 -197437
rect -96 -199631 -62 -198655
rect 62 -199631 96 -198655
rect -96 -200849 -62 -199873
rect 62 -200849 96 -199873
rect -96 -202067 -62 -201091
rect 62 -202067 96 -201091
rect -96 -203285 -62 -202309
rect 62 -203285 96 -202309
rect -96 -204503 -62 -203527
rect 62 -204503 96 -203527
rect -96 -205721 -62 -204745
rect 62 -205721 96 -204745
rect -96 -206939 -62 -205963
rect 62 -206939 96 -205963
rect -96 -208157 -62 -207181
rect 62 -208157 96 -207181
rect -96 -209375 -62 -208399
rect 62 -209375 96 -208399
rect -96 -210593 -62 -209617
rect 62 -210593 96 -209617
rect -96 -211811 -62 -210835
rect 62 -211811 96 -210835
rect -96 -213029 -62 -212053
rect 62 -213029 96 -212053
rect -96 -214247 -62 -213271
rect 62 -214247 96 -213271
rect -96 -215465 -62 -214489
rect 62 -215465 96 -214489
rect -96 -216683 -62 -215707
rect 62 -216683 96 -215707
rect -96 -217901 -62 -216925
rect 62 -217901 96 -216925
rect -96 -219119 -62 -218143
rect 62 -219119 96 -218143
rect -96 -220337 -62 -219361
rect 62 -220337 96 -219361
rect -96 -221555 -62 -220579
rect 62 -221555 96 -220579
rect -96 -222773 -62 -221797
rect 62 -222773 96 -221797
rect -96 -223991 -62 -223015
rect 62 -223991 96 -223015
rect -96 -225209 -62 -224233
rect 62 -225209 96 -224233
rect -96 -226427 -62 -225451
rect 62 -226427 96 -225451
rect -96 -227645 -62 -226669
rect 62 -227645 96 -226669
rect -96 -228863 -62 -227887
rect 62 -228863 96 -227887
rect -96 -230081 -62 -229105
rect 62 -230081 96 -229105
rect -96 -231299 -62 -230323
rect 62 -231299 96 -230323
rect -96 -232517 -62 -231541
rect 62 -232517 96 -231541
rect -96 -233735 -62 -232759
rect 62 -233735 96 -232759
rect -96 -234953 -62 -233977
rect 62 -234953 96 -233977
rect -96 -236171 -62 -235195
rect 62 -236171 96 -235195
rect -96 -237389 -62 -236413
rect 62 -237389 96 -236413
rect -96 -238607 -62 -237631
rect 62 -238607 96 -237631
rect -96 -239825 -62 -238849
rect 62 -239825 96 -238849
rect -96 -241043 -62 -240067
rect 62 -241043 96 -240067
rect -96 -242261 -62 -241285
rect 62 -242261 96 -241285
rect -96 -243479 -62 -242503
rect 62 -243479 96 -242503
rect -96 -244697 -62 -243721
rect 62 -244697 96 -243721
rect -96 -245915 -62 -244939
rect 62 -245915 96 -244939
rect -96 -247133 -62 -246157
rect 62 -247133 96 -246157
rect -96 -248351 -62 -247375
rect 62 -248351 96 -247375
rect -96 -249569 -62 -248593
rect 62 -249569 96 -248593
rect -96 -250787 -62 -249811
rect 62 -250787 96 -249811
rect -96 -252005 -62 -251029
rect 62 -252005 96 -251029
rect -96 -253223 -62 -252247
rect 62 -253223 96 -252247
rect -96 -254441 -62 -253465
rect 62 -254441 96 -253465
rect -96 -255659 -62 -254683
rect 62 -255659 96 -254683
rect -96 -256877 -62 -255901
rect 62 -256877 96 -255901
rect -96 -258095 -62 -257119
rect 62 -258095 96 -257119
rect -96 -259313 -62 -258337
rect 62 -259313 96 -258337
rect -96 -260531 -62 -259555
rect 62 -260531 96 -259555
rect -96 -261749 -62 -260773
rect 62 -261749 96 -260773
rect -96 -262967 -62 -261991
rect 62 -262967 96 -261991
rect -96 -264185 -62 -263209
rect 62 -264185 96 -263209
rect -96 -265403 -62 -264427
rect 62 -265403 96 -264427
rect -96 -266621 -62 -265645
rect 62 -266621 96 -265645
rect -96 -267839 -62 -266863
rect 62 -267839 96 -266863
rect -96 -269057 -62 -268081
rect 62 -269057 96 -268081
rect -96 -270275 -62 -269299
rect 62 -270275 96 -269299
rect -96 -271493 -62 -270517
rect 62 -271493 96 -270517
rect -96 -272711 -62 -271735
rect 62 -272711 96 -271735
rect -96 -273929 -62 -272953
rect 62 -273929 96 -272953
rect -96 -275147 -62 -274171
rect 62 -275147 96 -274171
rect -96 -276365 -62 -275389
rect 62 -276365 96 -275389
rect -96 -277583 -62 -276607
rect 62 -277583 96 -276607
rect -96 -278801 -62 -277825
rect 62 -278801 96 -277825
rect -96 -280019 -62 -279043
rect 62 -280019 96 -279043
rect -96 -281237 -62 -280261
rect 62 -281237 96 -280261
rect -96 -282455 -62 -281479
rect 62 -282455 96 -281479
rect -96 -283673 -62 -282697
rect 62 -283673 96 -282697
rect -96 -284891 -62 -283915
rect 62 -284891 96 -283915
rect -96 -286109 -62 -285133
rect 62 -286109 96 -285133
rect -96 -287327 -62 -286351
rect 62 -287327 96 -286351
rect -96 -288545 -62 -287569
rect 62 -288545 96 -287569
rect -96 -289763 -62 -288787
rect 62 -289763 96 -288787
rect -96 -290981 -62 -290005
rect 62 -290981 96 -290005
rect -96 -292199 -62 -291223
rect 62 -292199 96 -291223
rect -96 -293417 -62 -292441
rect 62 -293417 96 -292441
rect -96 -294635 -62 -293659
rect 62 -294635 96 -293659
rect -96 -295853 -62 -294877
rect 62 -295853 96 -294877
rect -96 -297071 -62 -296095
rect 62 -297071 96 -296095
rect -96 -298289 -62 -297313
rect 62 -298289 96 -297313
rect -96 -299507 -62 -298531
rect 62 -299507 96 -298531
rect -96 -300725 -62 -299749
rect 62 -300725 96 -299749
rect -96 -301943 -62 -300967
rect 62 -301943 96 -300967
rect -96 -303161 -62 -302185
rect 62 -303161 96 -302185
rect -96 -304379 -62 -303403
rect 62 -304379 96 -303403
rect -96 -305597 -62 -304621
rect 62 -305597 96 -304621
rect -96 -306815 -62 -305839
rect 62 -306815 96 -305839
rect -96 -308033 -62 -307057
rect 62 -308033 96 -307057
rect -96 -309251 -62 -308275
rect 62 -309251 96 -308275
rect -96 -310469 -62 -309493
rect 62 -310469 96 -309493
rect -96 -311687 -62 -310711
rect 62 -311687 96 -310711
rect -96 -312905 -62 -311929
rect 62 -312905 96 -311929
rect -96 -314123 -62 -313147
rect 62 -314123 96 -313147
rect -96 -315341 -62 -314365
rect 62 -315341 96 -314365
rect -96 -316559 -62 -315583
rect 62 -316559 96 -315583
rect -96 -317777 -62 -316801
rect 62 -317777 96 -316801
rect -96 -318995 -62 -318019
rect 62 -318995 96 -318019
rect -96 -320213 -62 -319237
rect 62 -320213 96 -319237
rect -96 -321431 -62 -320455
rect 62 -321431 96 -320455
rect -96 -322649 -62 -321673
rect 62 -322649 96 -321673
rect -96 -323867 -62 -322891
rect 62 -323867 96 -322891
rect -96 -325085 -62 -324109
rect 62 -325085 96 -324109
rect -96 -326303 -62 -325327
rect 62 -326303 96 -325327
rect -96 -327521 -62 -326545
rect 62 -327521 96 -326545
rect -96 -328739 -62 -327763
rect 62 -328739 96 -327763
rect -96 -329957 -62 -328981
rect 62 -329957 96 -328981
rect -96 -331175 -62 -330199
rect 62 -331175 96 -330199
rect -96 -332393 -62 -331417
rect 62 -332393 96 -331417
rect -96 -333611 -62 -332635
rect 62 -333611 96 -332635
rect -96 -334829 -62 -333853
rect 62 -334829 96 -333853
rect -96 -336047 -62 -335071
rect 62 -336047 96 -335071
rect -96 -337265 -62 -336289
rect 62 -337265 96 -336289
rect -96 -338483 -62 -337507
rect 62 -338483 96 -337507
rect -96 -339701 -62 -338725
rect 62 -339701 96 -338725
rect -96 -340919 -62 -339943
rect 62 -340919 96 -339943
rect -96 -342137 -62 -341161
rect 62 -342137 96 -341161
rect -96 -343355 -62 -342379
rect 62 -343355 96 -342379
rect -96 -344573 -62 -343597
rect 62 -344573 96 -343597
rect -96 -345791 -62 -344815
rect 62 -345791 96 -344815
rect -96 -347009 -62 -346033
rect 62 -347009 96 -346033
rect -96 -348227 -62 -347251
rect 62 -348227 96 -347251
rect -96 -349445 -62 -348469
rect 62 -349445 96 -348469
rect -96 -350663 -62 -349687
rect 62 -350663 96 -349687
rect -96 -351881 -62 -350905
rect 62 -351881 96 -350905
rect -96 -353099 -62 -352123
rect 62 -353099 96 -352123
rect -96 -354317 -62 -353341
rect 62 -354317 96 -353341
rect -96 -355535 -62 -354559
rect 62 -355535 96 -354559
rect -96 -356753 -62 -355777
rect 62 -356753 96 -355777
rect -96 -357971 -62 -356995
rect 62 -357971 96 -356995
rect -96 -359189 -62 -358213
rect 62 -359189 96 -358213
rect -96 -360407 -62 -359431
rect 62 -360407 96 -359431
rect -96 -361625 -62 -360649
rect 62 -361625 96 -360649
rect -96 -362843 -62 -361867
rect 62 -362843 96 -361867
rect -96 -364061 -62 -363085
rect 62 -364061 96 -363085
rect -96 -365279 -62 -364303
rect 62 -365279 96 -364303
rect -96 -366497 -62 -365521
rect 62 -366497 96 -365521
rect -96 -367715 -62 -366739
rect 62 -367715 96 -366739
rect -96 -368933 -62 -367957
rect 62 -368933 96 -367957
rect -96 -370151 -62 -369175
rect 62 -370151 96 -369175
rect -96 -371369 -62 -370393
rect 62 -371369 96 -370393
rect -96 -372587 -62 -371611
rect 62 -372587 96 -371611
rect -96 -373805 -62 -372829
rect 62 -373805 96 -372829
rect -96 -375023 -62 -374047
rect 62 -375023 96 -374047
rect -96 -376241 -62 -375265
rect 62 -376241 96 -375265
rect -96 -377459 -62 -376483
rect 62 -377459 96 -376483
rect -96 -378677 -62 -377701
rect 62 -378677 96 -377701
rect -96 -379895 -62 -378919
rect 62 -379895 96 -378919
rect -96 -381113 -62 -380137
rect 62 -381113 96 -380137
rect -96 -382331 -62 -381355
rect 62 -382331 96 -381355
rect -96 -383549 -62 -382573
rect 62 -383549 96 -382573
rect -96 -384767 -62 -383791
rect 62 -384767 96 -383791
rect -96 -385985 -62 -385009
rect 62 -385985 96 -385009
rect -96 -387203 -62 -386227
rect 62 -387203 96 -386227
rect -96 -388421 -62 -387445
rect 62 -388421 96 -387445
rect -96 -389639 -62 -388663
rect 62 -389639 96 -388663
rect -96 -390857 -62 -389881
rect 62 -390857 96 -389881
rect -96 -392075 -62 -391099
rect 62 -392075 96 -391099
rect -96 -393293 -62 -392317
rect 62 -393293 96 -392317
rect -96 -394511 -62 -393535
rect 62 -394511 96 -393535
rect -96 -395729 -62 -394753
rect 62 -395729 96 -394753
rect -96 -396947 -62 -395971
rect 62 -396947 96 -395971
rect -96 -398165 -62 -397189
rect 62 -398165 96 -397189
rect -96 -399383 -62 -398407
rect 62 -399383 96 -398407
rect -96 -400601 -62 -399625
rect 62 -400601 96 -399625
rect -96 -401819 -62 -400843
rect 62 -401819 96 -400843
rect -96 -403037 -62 -402061
rect 62 -403037 96 -402061
rect -96 -404255 -62 -403279
rect 62 -404255 96 -403279
rect -96 -405473 -62 -404497
rect 62 -405473 96 -404497
rect -96 -406691 -62 -405715
rect 62 -406691 96 -405715
rect -96 -407909 -62 -406933
rect 62 -407909 96 -406933
rect -96 -409127 -62 -408151
rect 62 -409127 96 -408151
rect -96 -410345 -62 -409369
rect 62 -410345 96 -409369
rect -96 -411563 -62 -410587
rect 62 -411563 96 -410587
rect -96 -412781 -62 -411805
rect 62 -412781 96 -411805
rect -96 -413999 -62 -413023
rect 62 -413999 96 -413023
rect -96 -415217 -62 -414241
rect 62 -415217 96 -414241
rect -96 -416435 -62 -415459
rect 62 -416435 96 -415459
rect -96 -417653 -62 -416677
rect 62 -417653 96 -416677
rect -96 -418871 -62 -417895
rect 62 -418871 96 -417895
rect -96 -420089 -62 -419113
rect 62 -420089 96 -419113
rect -96 -421307 -62 -420331
rect 62 -421307 96 -420331
rect -96 -422525 -62 -421549
rect 62 -422525 96 -421549
rect -96 -423743 -62 -422767
rect 62 -423743 96 -422767
rect -96 -424961 -62 -423985
rect 62 -424961 96 -423985
rect -96 -426179 -62 -425203
rect 62 -426179 96 -425203
rect -96 -427397 -62 -426421
rect 62 -427397 96 -426421
rect -96 -428615 -62 -427639
rect 62 -428615 96 -427639
rect -96 -429833 -62 -428857
rect 62 -429833 96 -428857
rect -96 -431051 -62 -430075
rect 62 -431051 96 -430075
rect -96 -432269 -62 -431293
rect 62 -432269 96 -431293
rect -96 -433487 -62 -432511
rect 62 -433487 96 -432511
rect -96 -434705 -62 -433729
rect 62 -434705 96 -433729
rect -96 -435923 -62 -434947
rect 62 -435923 96 -434947
rect -96 -437141 -62 -436165
rect 62 -437141 96 -436165
rect -96 -438359 -62 -437383
rect 62 -438359 96 -437383
rect -96 -439577 -62 -438601
rect 62 -439577 96 -438601
rect -96 -440795 -62 -439819
rect 62 -440795 96 -439819
rect -96 -442013 -62 -441037
rect 62 -442013 96 -441037
rect -96 -443231 -62 -442255
rect 62 -443231 96 -442255
rect -96 -444449 -62 -443473
rect 62 -444449 96 -443473
rect -96 -445667 -62 -444691
rect 62 -445667 96 -444691
rect -96 -446885 -62 -445909
rect 62 -446885 96 -445909
rect -96 -448103 -62 -447127
rect 62 -448103 96 -447127
rect -96 -449321 -62 -448345
rect 62 -449321 96 -448345
rect -96 -450539 -62 -449563
rect 62 -450539 96 -449563
rect -96 -451757 -62 -450781
rect 62 -451757 96 -450781
rect -96 -452975 -62 -451999
rect 62 -452975 96 -451999
rect -96 -454193 -62 -453217
rect 62 -454193 96 -453217
rect -96 -455411 -62 -454435
rect 62 -455411 96 -454435
rect -96 -456629 -62 -455653
rect 62 -456629 96 -455653
rect -96 -457847 -62 -456871
rect 62 -457847 96 -456871
rect -96 -459065 -62 -458089
rect 62 -459065 96 -458089
rect -96 -460283 -62 -459307
rect 62 -460283 96 -459307
rect -96 -461501 -62 -460525
rect 62 -461501 96 -460525
rect -96 -462719 -62 -461743
rect 62 -462719 96 -461743
rect -96 -463937 -62 -462961
rect 62 -463937 96 -462961
rect -96 -465155 -62 -464179
rect 62 -465155 96 -464179
rect -96 -466373 -62 -465397
rect 62 -466373 96 -465397
rect -96 -467591 -62 -466615
rect 62 -467591 96 -466615
rect -96 -468809 -62 -467833
rect 62 -468809 96 -467833
rect -96 -470027 -62 -469051
rect 62 -470027 96 -469051
rect -96 -471245 -62 -470269
rect 62 -471245 96 -470269
rect -96 -472463 -62 -471487
rect 62 -472463 96 -471487
rect -96 -473681 -62 -472705
rect 62 -473681 96 -472705
rect -96 -474899 -62 -473923
rect 62 -474899 96 -473923
rect -96 -476117 -62 -475141
rect 62 -476117 96 -475141
rect -96 -477335 -62 -476359
rect 62 -477335 96 -476359
rect -96 -478553 -62 -477577
rect 62 -478553 96 -477577
rect -96 -479771 -62 -478795
rect 62 -479771 96 -478795
rect -96 -480989 -62 -480013
rect 62 -480989 96 -480013
rect -96 -482207 -62 -481231
rect 62 -482207 96 -481231
rect -96 -483425 -62 -482449
rect 62 -483425 96 -482449
rect -96 -484643 -62 -483667
rect 62 -484643 96 -483667
rect -96 -485861 -62 -484885
rect 62 -485861 96 -484885
rect -96 -487079 -62 -486103
rect 62 -487079 96 -486103
rect -96 -488297 -62 -487321
rect 62 -488297 96 -487321
rect -96 -489515 -62 -488539
rect 62 -489515 96 -488539
rect -96 -490733 -62 -489757
rect 62 -490733 96 -489757
rect -96 -491951 -62 -490975
rect 62 -491951 96 -490975
rect -96 -493169 -62 -492193
rect 62 -493169 96 -492193
rect -96 -494387 -62 -493411
rect 62 -494387 96 -493411
rect -96 -495605 -62 -494629
rect 62 -495605 96 -494629
rect -96 -496823 -62 -495847
rect 62 -496823 96 -495847
rect -96 -498041 -62 -497065
rect 62 -498041 96 -497065
rect -96 -499259 -62 -498283
rect 62 -499259 96 -498283
rect -96 -500477 -62 -499501
rect 62 -500477 96 -499501
rect -96 -501695 -62 -500719
rect 62 -501695 96 -500719
rect -96 -502913 -62 -501937
rect 62 -502913 96 -501937
rect -96 -504131 -62 -503155
rect 62 -504131 96 -503155
rect -96 -505349 -62 -504373
rect 62 -505349 96 -504373
rect -96 -506567 -62 -505591
rect 62 -506567 96 -505591
rect -96 -507785 -62 -506809
rect 62 -507785 96 -506809
rect -96 -509003 -62 -508027
rect 62 -509003 96 -508027
rect -96 -510221 -62 -509245
rect 62 -510221 96 -509245
rect -96 -511439 -62 -510463
rect 62 -511439 96 -510463
rect -96 -512657 -62 -511681
rect 62 -512657 96 -511681
rect -96 -513875 -62 -512899
rect 62 -513875 96 -512899
rect -96 -515093 -62 -514117
rect 62 -515093 96 -514117
rect -96 -516311 -62 -515335
rect 62 -516311 96 -515335
rect -96 -517529 -62 -516553
rect 62 -517529 96 -516553
rect -96 -518747 -62 -517771
rect 62 -518747 96 -517771
rect -96 -519965 -62 -518989
rect 62 -519965 96 -518989
rect -96 -521183 -62 -520207
rect 62 -521183 96 -520207
rect -96 -522401 -62 -521425
rect 62 -522401 96 -521425
rect -96 -523619 -62 -522643
rect 62 -523619 96 -522643
rect -96 -524837 -62 -523861
rect 62 -524837 96 -523861
rect -96 -526055 -62 -525079
rect 62 -526055 96 -525079
rect -96 -527273 -62 -526297
rect 62 -527273 96 -526297
rect -96 -528491 -62 -527515
rect 62 -528491 96 -527515
rect -96 -529709 -62 -528733
rect 62 -529709 96 -528733
rect -96 -530927 -62 -529951
rect 62 -530927 96 -529951
rect -96 -532145 -62 -531169
rect 62 -532145 96 -531169
rect -96 -533363 -62 -532387
rect 62 -533363 96 -532387
rect -96 -534581 -62 -533605
rect 62 -534581 96 -533605
rect -96 -535799 -62 -534823
rect 62 -535799 96 -534823
rect -96 -537017 -62 -536041
rect 62 -537017 96 -536041
rect -96 -538235 -62 -537259
rect 62 -538235 96 -537259
rect -96 -539453 -62 -538477
rect 62 -539453 96 -538477
rect -96 -540671 -62 -539695
rect 62 -540671 96 -539695
rect -96 -541889 -62 -540913
rect 62 -541889 96 -540913
rect -96 -543107 -62 -542131
rect 62 -543107 96 -542131
rect -96 -544325 -62 -543349
rect 62 -544325 96 -543349
rect -96 -545543 -62 -544567
rect 62 -545543 96 -544567
rect -96 -546761 -62 -545785
rect 62 -546761 96 -545785
rect -96 -547979 -62 -547003
rect 62 -547979 96 -547003
rect -96 -549197 -62 -548221
rect 62 -549197 96 -548221
rect -96 -550415 -62 -549439
rect 62 -550415 96 -549439
rect -96 -551633 -62 -550657
rect 62 -551633 96 -550657
rect -96 -552851 -62 -551875
rect 62 -552851 96 -551875
rect -96 -554069 -62 -553093
rect 62 -554069 96 -553093
rect -96 -555287 -62 -554311
rect 62 -555287 96 -554311
rect -96 -556505 -62 -555529
rect 62 -556505 96 -555529
rect -96 -557723 -62 -556747
rect 62 -557723 96 -556747
rect -96 -558941 -62 -557965
rect 62 -558941 96 -557965
rect -96 -560159 -62 -559183
rect 62 -560159 96 -559183
rect -96 -561377 -62 -560401
rect 62 -561377 96 -560401
rect -96 -562595 -62 -561619
rect 62 -562595 96 -561619
rect -96 -563813 -62 -562837
rect 62 -563813 96 -562837
rect -96 -565031 -62 -564055
rect 62 -565031 96 -564055
rect -96 -566249 -62 -565273
rect 62 -566249 96 -565273
rect -96 -567467 -62 -566491
rect 62 -567467 96 -566491
rect -96 -568685 -62 -567709
rect 62 -568685 96 -567709
rect -96 -569903 -62 -568927
rect 62 -569903 96 -568927
rect -96 -571121 -62 -570145
rect 62 -571121 96 -570145
rect -96 -572339 -62 -571363
rect 62 -572339 96 -571363
rect -96 -573557 -62 -572581
rect 62 -573557 96 -572581
rect -96 -574775 -62 -573799
rect 62 -574775 96 -573799
rect -96 -575993 -62 -575017
rect 62 -575993 96 -575017
rect -96 -577211 -62 -576235
rect 62 -577211 96 -576235
rect -96 -578429 -62 -577453
rect 62 -578429 96 -577453
rect -96 -579647 -62 -578671
rect 62 -579647 96 -578671
rect -96 -580865 -62 -579889
rect 62 -580865 96 -579889
rect -96 -582083 -62 -581107
rect 62 -582083 96 -581107
rect -96 -583301 -62 -582325
rect 62 -583301 96 -582325
rect -96 -584519 -62 -583543
rect 62 -584519 96 -583543
rect -96 -585737 -62 -584761
rect 62 -585737 96 -584761
rect -96 -586955 -62 -585979
rect 62 -586955 96 -585979
rect -96 -588173 -62 -587197
rect 62 -588173 96 -587197
rect -96 -589391 -62 -588415
rect 62 -589391 96 -588415
rect -96 -590609 -62 -589633
rect 62 -590609 96 -589633
rect -96 -591827 -62 -590851
rect 62 -591827 96 -590851
rect -96 -593045 -62 -592069
rect 62 -593045 96 -592069
rect -96 -594263 -62 -593287
rect 62 -594263 96 -593287
rect -96 -595481 -62 -594505
rect 62 -595481 96 -594505
rect -96 -596699 -62 -595723
rect 62 -596699 96 -595723
rect -96 -597917 -62 -596941
rect 62 -597917 96 -596941
rect -96 -599135 -62 -598159
rect 62 -599135 96 -598159
rect -96 -600353 -62 -599377
rect 62 -600353 96 -599377
rect -96 -601571 -62 -600595
rect 62 -601571 96 -600595
rect -96 -602789 -62 -601813
rect 62 -602789 96 -601813
rect -96 -604007 -62 -603031
rect 62 -604007 96 -603031
rect -96 -605225 -62 -604249
rect 62 -605225 96 -604249
rect -96 -606443 -62 -605467
rect 62 -606443 96 -605467
rect -96 -607661 -62 -606685
rect 62 -607661 96 -606685
rect -96 -608879 -62 -607903
rect 62 -608879 96 -607903
<< mvpsubdiff >>
rect -242 609101 242 609113
rect -242 609067 -134 609101
rect 134 609067 242 609101
rect -242 609055 242 609067
rect -242 609005 -184 609055
rect -242 -609005 -230 609005
rect -196 -609005 -184 609005
rect 184 609005 242 609055
rect -242 -609055 -184 -609005
rect 184 -609005 196 609005
rect 230 -609005 242 609005
rect 184 -609055 242 -609005
rect -242 -609067 242 -609055
rect -242 -609101 -134 -609067
rect 134 -609101 242 -609067
rect -242 -609113 242 -609101
<< mvpsubdiffcont >>
rect -134 609067 134 609101
rect -230 -609005 -196 609005
rect 196 -609005 230 609005
rect -134 -609101 134 -609067
<< poly >>
rect -50 608963 50 608979
rect -50 608929 -34 608963
rect 34 608929 50 608963
rect -50 608891 50 608929
rect -50 607853 50 607891
rect -50 607819 -34 607853
rect 34 607819 50 607853
rect -50 607803 50 607819
rect -50 607745 50 607761
rect -50 607711 -34 607745
rect 34 607711 50 607745
rect -50 607673 50 607711
rect -50 606635 50 606673
rect -50 606601 -34 606635
rect 34 606601 50 606635
rect -50 606585 50 606601
rect -50 606527 50 606543
rect -50 606493 -34 606527
rect 34 606493 50 606527
rect -50 606455 50 606493
rect -50 605417 50 605455
rect -50 605383 -34 605417
rect 34 605383 50 605417
rect -50 605367 50 605383
rect -50 605309 50 605325
rect -50 605275 -34 605309
rect 34 605275 50 605309
rect -50 605237 50 605275
rect -50 604199 50 604237
rect -50 604165 -34 604199
rect 34 604165 50 604199
rect -50 604149 50 604165
rect -50 604091 50 604107
rect -50 604057 -34 604091
rect 34 604057 50 604091
rect -50 604019 50 604057
rect -50 602981 50 603019
rect -50 602947 -34 602981
rect 34 602947 50 602981
rect -50 602931 50 602947
rect -50 602873 50 602889
rect -50 602839 -34 602873
rect 34 602839 50 602873
rect -50 602801 50 602839
rect -50 601763 50 601801
rect -50 601729 -34 601763
rect 34 601729 50 601763
rect -50 601713 50 601729
rect -50 601655 50 601671
rect -50 601621 -34 601655
rect 34 601621 50 601655
rect -50 601583 50 601621
rect -50 600545 50 600583
rect -50 600511 -34 600545
rect 34 600511 50 600545
rect -50 600495 50 600511
rect -50 600437 50 600453
rect -50 600403 -34 600437
rect 34 600403 50 600437
rect -50 600365 50 600403
rect -50 599327 50 599365
rect -50 599293 -34 599327
rect 34 599293 50 599327
rect -50 599277 50 599293
rect -50 599219 50 599235
rect -50 599185 -34 599219
rect 34 599185 50 599219
rect -50 599147 50 599185
rect -50 598109 50 598147
rect -50 598075 -34 598109
rect 34 598075 50 598109
rect -50 598059 50 598075
rect -50 598001 50 598017
rect -50 597967 -34 598001
rect 34 597967 50 598001
rect -50 597929 50 597967
rect -50 596891 50 596929
rect -50 596857 -34 596891
rect 34 596857 50 596891
rect -50 596841 50 596857
rect -50 596783 50 596799
rect -50 596749 -34 596783
rect 34 596749 50 596783
rect -50 596711 50 596749
rect -50 595673 50 595711
rect -50 595639 -34 595673
rect 34 595639 50 595673
rect -50 595623 50 595639
rect -50 595565 50 595581
rect -50 595531 -34 595565
rect 34 595531 50 595565
rect -50 595493 50 595531
rect -50 594455 50 594493
rect -50 594421 -34 594455
rect 34 594421 50 594455
rect -50 594405 50 594421
rect -50 594347 50 594363
rect -50 594313 -34 594347
rect 34 594313 50 594347
rect -50 594275 50 594313
rect -50 593237 50 593275
rect -50 593203 -34 593237
rect 34 593203 50 593237
rect -50 593187 50 593203
rect -50 593129 50 593145
rect -50 593095 -34 593129
rect 34 593095 50 593129
rect -50 593057 50 593095
rect -50 592019 50 592057
rect -50 591985 -34 592019
rect 34 591985 50 592019
rect -50 591969 50 591985
rect -50 591911 50 591927
rect -50 591877 -34 591911
rect 34 591877 50 591911
rect -50 591839 50 591877
rect -50 590801 50 590839
rect -50 590767 -34 590801
rect 34 590767 50 590801
rect -50 590751 50 590767
rect -50 590693 50 590709
rect -50 590659 -34 590693
rect 34 590659 50 590693
rect -50 590621 50 590659
rect -50 589583 50 589621
rect -50 589549 -34 589583
rect 34 589549 50 589583
rect -50 589533 50 589549
rect -50 589475 50 589491
rect -50 589441 -34 589475
rect 34 589441 50 589475
rect -50 589403 50 589441
rect -50 588365 50 588403
rect -50 588331 -34 588365
rect 34 588331 50 588365
rect -50 588315 50 588331
rect -50 588257 50 588273
rect -50 588223 -34 588257
rect 34 588223 50 588257
rect -50 588185 50 588223
rect -50 587147 50 587185
rect -50 587113 -34 587147
rect 34 587113 50 587147
rect -50 587097 50 587113
rect -50 587039 50 587055
rect -50 587005 -34 587039
rect 34 587005 50 587039
rect -50 586967 50 587005
rect -50 585929 50 585967
rect -50 585895 -34 585929
rect 34 585895 50 585929
rect -50 585879 50 585895
rect -50 585821 50 585837
rect -50 585787 -34 585821
rect 34 585787 50 585821
rect -50 585749 50 585787
rect -50 584711 50 584749
rect -50 584677 -34 584711
rect 34 584677 50 584711
rect -50 584661 50 584677
rect -50 584603 50 584619
rect -50 584569 -34 584603
rect 34 584569 50 584603
rect -50 584531 50 584569
rect -50 583493 50 583531
rect -50 583459 -34 583493
rect 34 583459 50 583493
rect -50 583443 50 583459
rect -50 583385 50 583401
rect -50 583351 -34 583385
rect 34 583351 50 583385
rect -50 583313 50 583351
rect -50 582275 50 582313
rect -50 582241 -34 582275
rect 34 582241 50 582275
rect -50 582225 50 582241
rect -50 582167 50 582183
rect -50 582133 -34 582167
rect 34 582133 50 582167
rect -50 582095 50 582133
rect -50 581057 50 581095
rect -50 581023 -34 581057
rect 34 581023 50 581057
rect -50 581007 50 581023
rect -50 580949 50 580965
rect -50 580915 -34 580949
rect 34 580915 50 580949
rect -50 580877 50 580915
rect -50 579839 50 579877
rect -50 579805 -34 579839
rect 34 579805 50 579839
rect -50 579789 50 579805
rect -50 579731 50 579747
rect -50 579697 -34 579731
rect 34 579697 50 579731
rect -50 579659 50 579697
rect -50 578621 50 578659
rect -50 578587 -34 578621
rect 34 578587 50 578621
rect -50 578571 50 578587
rect -50 578513 50 578529
rect -50 578479 -34 578513
rect 34 578479 50 578513
rect -50 578441 50 578479
rect -50 577403 50 577441
rect -50 577369 -34 577403
rect 34 577369 50 577403
rect -50 577353 50 577369
rect -50 577295 50 577311
rect -50 577261 -34 577295
rect 34 577261 50 577295
rect -50 577223 50 577261
rect -50 576185 50 576223
rect -50 576151 -34 576185
rect 34 576151 50 576185
rect -50 576135 50 576151
rect -50 576077 50 576093
rect -50 576043 -34 576077
rect 34 576043 50 576077
rect -50 576005 50 576043
rect -50 574967 50 575005
rect -50 574933 -34 574967
rect 34 574933 50 574967
rect -50 574917 50 574933
rect -50 574859 50 574875
rect -50 574825 -34 574859
rect 34 574825 50 574859
rect -50 574787 50 574825
rect -50 573749 50 573787
rect -50 573715 -34 573749
rect 34 573715 50 573749
rect -50 573699 50 573715
rect -50 573641 50 573657
rect -50 573607 -34 573641
rect 34 573607 50 573641
rect -50 573569 50 573607
rect -50 572531 50 572569
rect -50 572497 -34 572531
rect 34 572497 50 572531
rect -50 572481 50 572497
rect -50 572423 50 572439
rect -50 572389 -34 572423
rect 34 572389 50 572423
rect -50 572351 50 572389
rect -50 571313 50 571351
rect -50 571279 -34 571313
rect 34 571279 50 571313
rect -50 571263 50 571279
rect -50 571205 50 571221
rect -50 571171 -34 571205
rect 34 571171 50 571205
rect -50 571133 50 571171
rect -50 570095 50 570133
rect -50 570061 -34 570095
rect 34 570061 50 570095
rect -50 570045 50 570061
rect -50 569987 50 570003
rect -50 569953 -34 569987
rect 34 569953 50 569987
rect -50 569915 50 569953
rect -50 568877 50 568915
rect -50 568843 -34 568877
rect 34 568843 50 568877
rect -50 568827 50 568843
rect -50 568769 50 568785
rect -50 568735 -34 568769
rect 34 568735 50 568769
rect -50 568697 50 568735
rect -50 567659 50 567697
rect -50 567625 -34 567659
rect 34 567625 50 567659
rect -50 567609 50 567625
rect -50 567551 50 567567
rect -50 567517 -34 567551
rect 34 567517 50 567551
rect -50 567479 50 567517
rect -50 566441 50 566479
rect -50 566407 -34 566441
rect 34 566407 50 566441
rect -50 566391 50 566407
rect -50 566333 50 566349
rect -50 566299 -34 566333
rect 34 566299 50 566333
rect -50 566261 50 566299
rect -50 565223 50 565261
rect -50 565189 -34 565223
rect 34 565189 50 565223
rect -50 565173 50 565189
rect -50 565115 50 565131
rect -50 565081 -34 565115
rect 34 565081 50 565115
rect -50 565043 50 565081
rect -50 564005 50 564043
rect -50 563971 -34 564005
rect 34 563971 50 564005
rect -50 563955 50 563971
rect -50 563897 50 563913
rect -50 563863 -34 563897
rect 34 563863 50 563897
rect -50 563825 50 563863
rect -50 562787 50 562825
rect -50 562753 -34 562787
rect 34 562753 50 562787
rect -50 562737 50 562753
rect -50 562679 50 562695
rect -50 562645 -34 562679
rect 34 562645 50 562679
rect -50 562607 50 562645
rect -50 561569 50 561607
rect -50 561535 -34 561569
rect 34 561535 50 561569
rect -50 561519 50 561535
rect -50 561461 50 561477
rect -50 561427 -34 561461
rect 34 561427 50 561461
rect -50 561389 50 561427
rect -50 560351 50 560389
rect -50 560317 -34 560351
rect 34 560317 50 560351
rect -50 560301 50 560317
rect -50 560243 50 560259
rect -50 560209 -34 560243
rect 34 560209 50 560243
rect -50 560171 50 560209
rect -50 559133 50 559171
rect -50 559099 -34 559133
rect 34 559099 50 559133
rect -50 559083 50 559099
rect -50 559025 50 559041
rect -50 558991 -34 559025
rect 34 558991 50 559025
rect -50 558953 50 558991
rect -50 557915 50 557953
rect -50 557881 -34 557915
rect 34 557881 50 557915
rect -50 557865 50 557881
rect -50 557807 50 557823
rect -50 557773 -34 557807
rect 34 557773 50 557807
rect -50 557735 50 557773
rect -50 556697 50 556735
rect -50 556663 -34 556697
rect 34 556663 50 556697
rect -50 556647 50 556663
rect -50 556589 50 556605
rect -50 556555 -34 556589
rect 34 556555 50 556589
rect -50 556517 50 556555
rect -50 555479 50 555517
rect -50 555445 -34 555479
rect 34 555445 50 555479
rect -50 555429 50 555445
rect -50 555371 50 555387
rect -50 555337 -34 555371
rect 34 555337 50 555371
rect -50 555299 50 555337
rect -50 554261 50 554299
rect -50 554227 -34 554261
rect 34 554227 50 554261
rect -50 554211 50 554227
rect -50 554153 50 554169
rect -50 554119 -34 554153
rect 34 554119 50 554153
rect -50 554081 50 554119
rect -50 553043 50 553081
rect -50 553009 -34 553043
rect 34 553009 50 553043
rect -50 552993 50 553009
rect -50 552935 50 552951
rect -50 552901 -34 552935
rect 34 552901 50 552935
rect -50 552863 50 552901
rect -50 551825 50 551863
rect -50 551791 -34 551825
rect 34 551791 50 551825
rect -50 551775 50 551791
rect -50 551717 50 551733
rect -50 551683 -34 551717
rect 34 551683 50 551717
rect -50 551645 50 551683
rect -50 550607 50 550645
rect -50 550573 -34 550607
rect 34 550573 50 550607
rect -50 550557 50 550573
rect -50 550499 50 550515
rect -50 550465 -34 550499
rect 34 550465 50 550499
rect -50 550427 50 550465
rect -50 549389 50 549427
rect -50 549355 -34 549389
rect 34 549355 50 549389
rect -50 549339 50 549355
rect -50 549281 50 549297
rect -50 549247 -34 549281
rect 34 549247 50 549281
rect -50 549209 50 549247
rect -50 548171 50 548209
rect -50 548137 -34 548171
rect 34 548137 50 548171
rect -50 548121 50 548137
rect -50 548063 50 548079
rect -50 548029 -34 548063
rect 34 548029 50 548063
rect -50 547991 50 548029
rect -50 546953 50 546991
rect -50 546919 -34 546953
rect 34 546919 50 546953
rect -50 546903 50 546919
rect -50 546845 50 546861
rect -50 546811 -34 546845
rect 34 546811 50 546845
rect -50 546773 50 546811
rect -50 545735 50 545773
rect -50 545701 -34 545735
rect 34 545701 50 545735
rect -50 545685 50 545701
rect -50 545627 50 545643
rect -50 545593 -34 545627
rect 34 545593 50 545627
rect -50 545555 50 545593
rect -50 544517 50 544555
rect -50 544483 -34 544517
rect 34 544483 50 544517
rect -50 544467 50 544483
rect -50 544409 50 544425
rect -50 544375 -34 544409
rect 34 544375 50 544409
rect -50 544337 50 544375
rect -50 543299 50 543337
rect -50 543265 -34 543299
rect 34 543265 50 543299
rect -50 543249 50 543265
rect -50 543191 50 543207
rect -50 543157 -34 543191
rect 34 543157 50 543191
rect -50 543119 50 543157
rect -50 542081 50 542119
rect -50 542047 -34 542081
rect 34 542047 50 542081
rect -50 542031 50 542047
rect -50 541973 50 541989
rect -50 541939 -34 541973
rect 34 541939 50 541973
rect -50 541901 50 541939
rect -50 540863 50 540901
rect -50 540829 -34 540863
rect 34 540829 50 540863
rect -50 540813 50 540829
rect -50 540755 50 540771
rect -50 540721 -34 540755
rect 34 540721 50 540755
rect -50 540683 50 540721
rect -50 539645 50 539683
rect -50 539611 -34 539645
rect 34 539611 50 539645
rect -50 539595 50 539611
rect -50 539537 50 539553
rect -50 539503 -34 539537
rect 34 539503 50 539537
rect -50 539465 50 539503
rect -50 538427 50 538465
rect -50 538393 -34 538427
rect 34 538393 50 538427
rect -50 538377 50 538393
rect -50 538319 50 538335
rect -50 538285 -34 538319
rect 34 538285 50 538319
rect -50 538247 50 538285
rect -50 537209 50 537247
rect -50 537175 -34 537209
rect 34 537175 50 537209
rect -50 537159 50 537175
rect -50 537101 50 537117
rect -50 537067 -34 537101
rect 34 537067 50 537101
rect -50 537029 50 537067
rect -50 535991 50 536029
rect -50 535957 -34 535991
rect 34 535957 50 535991
rect -50 535941 50 535957
rect -50 535883 50 535899
rect -50 535849 -34 535883
rect 34 535849 50 535883
rect -50 535811 50 535849
rect -50 534773 50 534811
rect -50 534739 -34 534773
rect 34 534739 50 534773
rect -50 534723 50 534739
rect -50 534665 50 534681
rect -50 534631 -34 534665
rect 34 534631 50 534665
rect -50 534593 50 534631
rect -50 533555 50 533593
rect -50 533521 -34 533555
rect 34 533521 50 533555
rect -50 533505 50 533521
rect -50 533447 50 533463
rect -50 533413 -34 533447
rect 34 533413 50 533447
rect -50 533375 50 533413
rect -50 532337 50 532375
rect -50 532303 -34 532337
rect 34 532303 50 532337
rect -50 532287 50 532303
rect -50 532229 50 532245
rect -50 532195 -34 532229
rect 34 532195 50 532229
rect -50 532157 50 532195
rect -50 531119 50 531157
rect -50 531085 -34 531119
rect 34 531085 50 531119
rect -50 531069 50 531085
rect -50 531011 50 531027
rect -50 530977 -34 531011
rect 34 530977 50 531011
rect -50 530939 50 530977
rect -50 529901 50 529939
rect -50 529867 -34 529901
rect 34 529867 50 529901
rect -50 529851 50 529867
rect -50 529793 50 529809
rect -50 529759 -34 529793
rect 34 529759 50 529793
rect -50 529721 50 529759
rect -50 528683 50 528721
rect -50 528649 -34 528683
rect 34 528649 50 528683
rect -50 528633 50 528649
rect -50 528575 50 528591
rect -50 528541 -34 528575
rect 34 528541 50 528575
rect -50 528503 50 528541
rect -50 527465 50 527503
rect -50 527431 -34 527465
rect 34 527431 50 527465
rect -50 527415 50 527431
rect -50 527357 50 527373
rect -50 527323 -34 527357
rect 34 527323 50 527357
rect -50 527285 50 527323
rect -50 526247 50 526285
rect -50 526213 -34 526247
rect 34 526213 50 526247
rect -50 526197 50 526213
rect -50 526139 50 526155
rect -50 526105 -34 526139
rect 34 526105 50 526139
rect -50 526067 50 526105
rect -50 525029 50 525067
rect -50 524995 -34 525029
rect 34 524995 50 525029
rect -50 524979 50 524995
rect -50 524921 50 524937
rect -50 524887 -34 524921
rect 34 524887 50 524921
rect -50 524849 50 524887
rect -50 523811 50 523849
rect -50 523777 -34 523811
rect 34 523777 50 523811
rect -50 523761 50 523777
rect -50 523703 50 523719
rect -50 523669 -34 523703
rect 34 523669 50 523703
rect -50 523631 50 523669
rect -50 522593 50 522631
rect -50 522559 -34 522593
rect 34 522559 50 522593
rect -50 522543 50 522559
rect -50 522485 50 522501
rect -50 522451 -34 522485
rect 34 522451 50 522485
rect -50 522413 50 522451
rect -50 521375 50 521413
rect -50 521341 -34 521375
rect 34 521341 50 521375
rect -50 521325 50 521341
rect -50 521267 50 521283
rect -50 521233 -34 521267
rect 34 521233 50 521267
rect -50 521195 50 521233
rect -50 520157 50 520195
rect -50 520123 -34 520157
rect 34 520123 50 520157
rect -50 520107 50 520123
rect -50 520049 50 520065
rect -50 520015 -34 520049
rect 34 520015 50 520049
rect -50 519977 50 520015
rect -50 518939 50 518977
rect -50 518905 -34 518939
rect 34 518905 50 518939
rect -50 518889 50 518905
rect -50 518831 50 518847
rect -50 518797 -34 518831
rect 34 518797 50 518831
rect -50 518759 50 518797
rect -50 517721 50 517759
rect -50 517687 -34 517721
rect 34 517687 50 517721
rect -50 517671 50 517687
rect -50 517613 50 517629
rect -50 517579 -34 517613
rect 34 517579 50 517613
rect -50 517541 50 517579
rect -50 516503 50 516541
rect -50 516469 -34 516503
rect 34 516469 50 516503
rect -50 516453 50 516469
rect -50 516395 50 516411
rect -50 516361 -34 516395
rect 34 516361 50 516395
rect -50 516323 50 516361
rect -50 515285 50 515323
rect -50 515251 -34 515285
rect 34 515251 50 515285
rect -50 515235 50 515251
rect -50 515177 50 515193
rect -50 515143 -34 515177
rect 34 515143 50 515177
rect -50 515105 50 515143
rect -50 514067 50 514105
rect -50 514033 -34 514067
rect 34 514033 50 514067
rect -50 514017 50 514033
rect -50 513959 50 513975
rect -50 513925 -34 513959
rect 34 513925 50 513959
rect -50 513887 50 513925
rect -50 512849 50 512887
rect -50 512815 -34 512849
rect 34 512815 50 512849
rect -50 512799 50 512815
rect -50 512741 50 512757
rect -50 512707 -34 512741
rect 34 512707 50 512741
rect -50 512669 50 512707
rect -50 511631 50 511669
rect -50 511597 -34 511631
rect 34 511597 50 511631
rect -50 511581 50 511597
rect -50 511523 50 511539
rect -50 511489 -34 511523
rect 34 511489 50 511523
rect -50 511451 50 511489
rect -50 510413 50 510451
rect -50 510379 -34 510413
rect 34 510379 50 510413
rect -50 510363 50 510379
rect -50 510305 50 510321
rect -50 510271 -34 510305
rect 34 510271 50 510305
rect -50 510233 50 510271
rect -50 509195 50 509233
rect -50 509161 -34 509195
rect 34 509161 50 509195
rect -50 509145 50 509161
rect -50 509087 50 509103
rect -50 509053 -34 509087
rect 34 509053 50 509087
rect -50 509015 50 509053
rect -50 507977 50 508015
rect -50 507943 -34 507977
rect 34 507943 50 507977
rect -50 507927 50 507943
rect -50 507869 50 507885
rect -50 507835 -34 507869
rect 34 507835 50 507869
rect -50 507797 50 507835
rect -50 506759 50 506797
rect -50 506725 -34 506759
rect 34 506725 50 506759
rect -50 506709 50 506725
rect -50 506651 50 506667
rect -50 506617 -34 506651
rect 34 506617 50 506651
rect -50 506579 50 506617
rect -50 505541 50 505579
rect -50 505507 -34 505541
rect 34 505507 50 505541
rect -50 505491 50 505507
rect -50 505433 50 505449
rect -50 505399 -34 505433
rect 34 505399 50 505433
rect -50 505361 50 505399
rect -50 504323 50 504361
rect -50 504289 -34 504323
rect 34 504289 50 504323
rect -50 504273 50 504289
rect -50 504215 50 504231
rect -50 504181 -34 504215
rect 34 504181 50 504215
rect -50 504143 50 504181
rect -50 503105 50 503143
rect -50 503071 -34 503105
rect 34 503071 50 503105
rect -50 503055 50 503071
rect -50 502997 50 503013
rect -50 502963 -34 502997
rect 34 502963 50 502997
rect -50 502925 50 502963
rect -50 501887 50 501925
rect -50 501853 -34 501887
rect 34 501853 50 501887
rect -50 501837 50 501853
rect -50 501779 50 501795
rect -50 501745 -34 501779
rect 34 501745 50 501779
rect -50 501707 50 501745
rect -50 500669 50 500707
rect -50 500635 -34 500669
rect 34 500635 50 500669
rect -50 500619 50 500635
rect -50 500561 50 500577
rect -50 500527 -34 500561
rect 34 500527 50 500561
rect -50 500489 50 500527
rect -50 499451 50 499489
rect -50 499417 -34 499451
rect 34 499417 50 499451
rect -50 499401 50 499417
rect -50 499343 50 499359
rect -50 499309 -34 499343
rect 34 499309 50 499343
rect -50 499271 50 499309
rect -50 498233 50 498271
rect -50 498199 -34 498233
rect 34 498199 50 498233
rect -50 498183 50 498199
rect -50 498125 50 498141
rect -50 498091 -34 498125
rect 34 498091 50 498125
rect -50 498053 50 498091
rect -50 497015 50 497053
rect -50 496981 -34 497015
rect 34 496981 50 497015
rect -50 496965 50 496981
rect -50 496907 50 496923
rect -50 496873 -34 496907
rect 34 496873 50 496907
rect -50 496835 50 496873
rect -50 495797 50 495835
rect -50 495763 -34 495797
rect 34 495763 50 495797
rect -50 495747 50 495763
rect -50 495689 50 495705
rect -50 495655 -34 495689
rect 34 495655 50 495689
rect -50 495617 50 495655
rect -50 494579 50 494617
rect -50 494545 -34 494579
rect 34 494545 50 494579
rect -50 494529 50 494545
rect -50 494471 50 494487
rect -50 494437 -34 494471
rect 34 494437 50 494471
rect -50 494399 50 494437
rect -50 493361 50 493399
rect -50 493327 -34 493361
rect 34 493327 50 493361
rect -50 493311 50 493327
rect -50 493253 50 493269
rect -50 493219 -34 493253
rect 34 493219 50 493253
rect -50 493181 50 493219
rect -50 492143 50 492181
rect -50 492109 -34 492143
rect 34 492109 50 492143
rect -50 492093 50 492109
rect -50 492035 50 492051
rect -50 492001 -34 492035
rect 34 492001 50 492035
rect -50 491963 50 492001
rect -50 490925 50 490963
rect -50 490891 -34 490925
rect 34 490891 50 490925
rect -50 490875 50 490891
rect -50 490817 50 490833
rect -50 490783 -34 490817
rect 34 490783 50 490817
rect -50 490745 50 490783
rect -50 489707 50 489745
rect -50 489673 -34 489707
rect 34 489673 50 489707
rect -50 489657 50 489673
rect -50 489599 50 489615
rect -50 489565 -34 489599
rect 34 489565 50 489599
rect -50 489527 50 489565
rect -50 488489 50 488527
rect -50 488455 -34 488489
rect 34 488455 50 488489
rect -50 488439 50 488455
rect -50 488381 50 488397
rect -50 488347 -34 488381
rect 34 488347 50 488381
rect -50 488309 50 488347
rect -50 487271 50 487309
rect -50 487237 -34 487271
rect 34 487237 50 487271
rect -50 487221 50 487237
rect -50 487163 50 487179
rect -50 487129 -34 487163
rect 34 487129 50 487163
rect -50 487091 50 487129
rect -50 486053 50 486091
rect -50 486019 -34 486053
rect 34 486019 50 486053
rect -50 486003 50 486019
rect -50 485945 50 485961
rect -50 485911 -34 485945
rect 34 485911 50 485945
rect -50 485873 50 485911
rect -50 484835 50 484873
rect -50 484801 -34 484835
rect 34 484801 50 484835
rect -50 484785 50 484801
rect -50 484727 50 484743
rect -50 484693 -34 484727
rect 34 484693 50 484727
rect -50 484655 50 484693
rect -50 483617 50 483655
rect -50 483583 -34 483617
rect 34 483583 50 483617
rect -50 483567 50 483583
rect -50 483509 50 483525
rect -50 483475 -34 483509
rect 34 483475 50 483509
rect -50 483437 50 483475
rect -50 482399 50 482437
rect -50 482365 -34 482399
rect 34 482365 50 482399
rect -50 482349 50 482365
rect -50 482291 50 482307
rect -50 482257 -34 482291
rect 34 482257 50 482291
rect -50 482219 50 482257
rect -50 481181 50 481219
rect -50 481147 -34 481181
rect 34 481147 50 481181
rect -50 481131 50 481147
rect -50 481073 50 481089
rect -50 481039 -34 481073
rect 34 481039 50 481073
rect -50 481001 50 481039
rect -50 479963 50 480001
rect -50 479929 -34 479963
rect 34 479929 50 479963
rect -50 479913 50 479929
rect -50 479855 50 479871
rect -50 479821 -34 479855
rect 34 479821 50 479855
rect -50 479783 50 479821
rect -50 478745 50 478783
rect -50 478711 -34 478745
rect 34 478711 50 478745
rect -50 478695 50 478711
rect -50 478637 50 478653
rect -50 478603 -34 478637
rect 34 478603 50 478637
rect -50 478565 50 478603
rect -50 477527 50 477565
rect -50 477493 -34 477527
rect 34 477493 50 477527
rect -50 477477 50 477493
rect -50 477419 50 477435
rect -50 477385 -34 477419
rect 34 477385 50 477419
rect -50 477347 50 477385
rect -50 476309 50 476347
rect -50 476275 -34 476309
rect 34 476275 50 476309
rect -50 476259 50 476275
rect -50 476201 50 476217
rect -50 476167 -34 476201
rect 34 476167 50 476201
rect -50 476129 50 476167
rect -50 475091 50 475129
rect -50 475057 -34 475091
rect 34 475057 50 475091
rect -50 475041 50 475057
rect -50 474983 50 474999
rect -50 474949 -34 474983
rect 34 474949 50 474983
rect -50 474911 50 474949
rect -50 473873 50 473911
rect -50 473839 -34 473873
rect 34 473839 50 473873
rect -50 473823 50 473839
rect -50 473765 50 473781
rect -50 473731 -34 473765
rect 34 473731 50 473765
rect -50 473693 50 473731
rect -50 472655 50 472693
rect -50 472621 -34 472655
rect 34 472621 50 472655
rect -50 472605 50 472621
rect -50 472547 50 472563
rect -50 472513 -34 472547
rect 34 472513 50 472547
rect -50 472475 50 472513
rect -50 471437 50 471475
rect -50 471403 -34 471437
rect 34 471403 50 471437
rect -50 471387 50 471403
rect -50 471329 50 471345
rect -50 471295 -34 471329
rect 34 471295 50 471329
rect -50 471257 50 471295
rect -50 470219 50 470257
rect -50 470185 -34 470219
rect 34 470185 50 470219
rect -50 470169 50 470185
rect -50 470111 50 470127
rect -50 470077 -34 470111
rect 34 470077 50 470111
rect -50 470039 50 470077
rect -50 469001 50 469039
rect -50 468967 -34 469001
rect 34 468967 50 469001
rect -50 468951 50 468967
rect -50 468893 50 468909
rect -50 468859 -34 468893
rect 34 468859 50 468893
rect -50 468821 50 468859
rect -50 467783 50 467821
rect -50 467749 -34 467783
rect 34 467749 50 467783
rect -50 467733 50 467749
rect -50 467675 50 467691
rect -50 467641 -34 467675
rect 34 467641 50 467675
rect -50 467603 50 467641
rect -50 466565 50 466603
rect -50 466531 -34 466565
rect 34 466531 50 466565
rect -50 466515 50 466531
rect -50 466457 50 466473
rect -50 466423 -34 466457
rect 34 466423 50 466457
rect -50 466385 50 466423
rect -50 465347 50 465385
rect -50 465313 -34 465347
rect 34 465313 50 465347
rect -50 465297 50 465313
rect -50 465239 50 465255
rect -50 465205 -34 465239
rect 34 465205 50 465239
rect -50 465167 50 465205
rect -50 464129 50 464167
rect -50 464095 -34 464129
rect 34 464095 50 464129
rect -50 464079 50 464095
rect -50 464021 50 464037
rect -50 463987 -34 464021
rect 34 463987 50 464021
rect -50 463949 50 463987
rect -50 462911 50 462949
rect -50 462877 -34 462911
rect 34 462877 50 462911
rect -50 462861 50 462877
rect -50 462803 50 462819
rect -50 462769 -34 462803
rect 34 462769 50 462803
rect -50 462731 50 462769
rect -50 461693 50 461731
rect -50 461659 -34 461693
rect 34 461659 50 461693
rect -50 461643 50 461659
rect -50 461585 50 461601
rect -50 461551 -34 461585
rect 34 461551 50 461585
rect -50 461513 50 461551
rect -50 460475 50 460513
rect -50 460441 -34 460475
rect 34 460441 50 460475
rect -50 460425 50 460441
rect -50 460367 50 460383
rect -50 460333 -34 460367
rect 34 460333 50 460367
rect -50 460295 50 460333
rect -50 459257 50 459295
rect -50 459223 -34 459257
rect 34 459223 50 459257
rect -50 459207 50 459223
rect -50 459149 50 459165
rect -50 459115 -34 459149
rect 34 459115 50 459149
rect -50 459077 50 459115
rect -50 458039 50 458077
rect -50 458005 -34 458039
rect 34 458005 50 458039
rect -50 457989 50 458005
rect -50 457931 50 457947
rect -50 457897 -34 457931
rect 34 457897 50 457931
rect -50 457859 50 457897
rect -50 456821 50 456859
rect -50 456787 -34 456821
rect 34 456787 50 456821
rect -50 456771 50 456787
rect -50 456713 50 456729
rect -50 456679 -34 456713
rect 34 456679 50 456713
rect -50 456641 50 456679
rect -50 455603 50 455641
rect -50 455569 -34 455603
rect 34 455569 50 455603
rect -50 455553 50 455569
rect -50 455495 50 455511
rect -50 455461 -34 455495
rect 34 455461 50 455495
rect -50 455423 50 455461
rect -50 454385 50 454423
rect -50 454351 -34 454385
rect 34 454351 50 454385
rect -50 454335 50 454351
rect -50 454277 50 454293
rect -50 454243 -34 454277
rect 34 454243 50 454277
rect -50 454205 50 454243
rect -50 453167 50 453205
rect -50 453133 -34 453167
rect 34 453133 50 453167
rect -50 453117 50 453133
rect -50 453059 50 453075
rect -50 453025 -34 453059
rect 34 453025 50 453059
rect -50 452987 50 453025
rect -50 451949 50 451987
rect -50 451915 -34 451949
rect 34 451915 50 451949
rect -50 451899 50 451915
rect -50 451841 50 451857
rect -50 451807 -34 451841
rect 34 451807 50 451841
rect -50 451769 50 451807
rect -50 450731 50 450769
rect -50 450697 -34 450731
rect 34 450697 50 450731
rect -50 450681 50 450697
rect -50 450623 50 450639
rect -50 450589 -34 450623
rect 34 450589 50 450623
rect -50 450551 50 450589
rect -50 449513 50 449551
rect -50 449479 -34 449513
rect 34 449479 50 449513
rect -50 449463 50 449479
rect -50 449405 50 449421
rect -50 449371 -34 449405
rect 34 449371 50 449405
rect -50 449333 50 449371
rect -50 448295 50 448333
rect -50 448261 -34 448295
rect 34 448261 50 448295
rect -50 448245 50 448261
rect -50 448187 50 448203
rect -50 448153 -34 448187
rect 34 448153 50 448187
rect -50 448115 50 448153
rect -50 447077 50 447115
rect -50 447043 -34 447077
rect 34 447043 50 447077
rect -50 447027 50 447043
rect -50 446969 50 446985
rect -50 446935 -34 446969
rect 34 446935 50 446969
rect -50 446897 50 446935
rect -50 445859 50 445897
rect -50 445825 -34 445859
rect 34 445825 50 445859
rect -50 445809 50 445825
rect -50 445751 50 445767
rect -50 445717 -34 445751
rect 34 445717 50 445751
rect -50 445679 50 445717
rect -50 444641 50 444679
rect -50 444607 -34 444641
rect 34 444607 50 444641
rect -50 444591 50 444607
rect -50 444533 50 444549
rect -50 444499 -34 444533
rect 34 444499 50 444533
rect -50 444461 50 444499
rect -50 443423 50 443461
rect -50 443389 -34 443423
rect 34 443389 50 443423
rect -50 443373 50 443389
rect -50 443315 50 443331
rect -50 443281 -34 443315
rect 34 443281 50 443315
rect -50 443243 50 443281
rect -50 442205 50 442243
rect -50 442171 -34 442205
rect 34 442171 50 442205
rect -50 442155 50 442171
rect -50 442097 50 442113
rect -50 442063 -34 442097
rect 34 442063 50 442097
rect -50 442025 50 442063
rect -50 440987 50 441025
rect -50 440953 -34 440987
rect 34 440953 50 440987
rect -50 440937 50 440953
rect -50 440879 50 440895
rect -50 440845 -34 440879
rect 34 440845 50 440879
rect -50 440807 50 440845
rect -50 439769 50 439807
rect -50 439735 -34 439769
rect 34 439735 50 439769
rect -50 439719 50 439735
rect -50 439661 50 439677
rect -50 439627 -34 439661
rect 34 439627 50 439661
rect -50 439589 50 439627
rect -50 438551 50 438589
rect -50 438517 -34 438551
rect 34 438517 50 438551
rect -50 438501 50 438517
rect -50 438443 50 438459
rect -50 438409 -34 438443
rect 34 438409 50 438443
rect -50 438371 50 438409
rect -50 437333 50 437371
rect -50 437299 -34 437333
rect 34 437299 50 437333
rect -50 437283 50 437299
rect -50 437225 50 437241
rect -50 437191 -34 437225
rect 34 437191 50 437225
rect -50 437153 50 437191
rect -50 436115 50 436153
rect -50 436081 -34 436115
rect 34 436081 50 436115
rect -50 436065 50 436081
rect -50 436007 50 436023
rect -50 435973 -34 436007
rect 34 435973 50 436007
rect -50 435935 50 435973
rect -50 434897 50 434935
rect -50 434863 -34 434897
rect 34 434863 50 434897
rect -50 434847 50 434863
rect -50 434789 50 434805
rect -50 434755 -34 434789
rect 34 434755 50 434789
rect -50 434717 50 434755
rect -50 433679 50 433717
rect -50 433645 -34 433679
rect 34 433645 50 433679
rect -50 433629 50 433645
rect -50 433571 50 433587
rect -50 433537 -34 433571
rect 34 433537 50 433571
rect -50 433499 50 433537
rect -50 432461 50 432499
rect -50 432427 -34 432461
rect 34 432427 50 432461
rect -50 432411 50 432427
rect -50 432353 50 432369
rect -50 432319 -34 432353
rect 34 432319 50 432353
rect -50 432281 50 432319
rect -50 431243 50 431281
rect -50 431209 -34 431243
rect 34 431209 50 431243
rect -50 431193 50 431209
rect -50 431135 50 431151
rect -50 431101 -34 431135
rect 34 431101 50 431135
rect -50 431063 50 431101
rect -50 430025 50 430063
rect -50 429991 -34 430025
rect 34 429991 50 430025
rect -50 429975 50 429991
rect -50 429917 50 429933
rect -50 429883 -34 429917
rect 34 429883 50 429917
rect -50 429845 50 429883
rect -50 428807 50 428845
rect -50 428773 -34 428807
rect 34 428773 50 428807
rect -50 428757 50 428773
rect -50 428699 50 428715
rect -50 428665 -34 428699
rect 34 428665 50 428699
rect -50 428627 50 428665
rect -50 427589 50 427627
rect -50 427555 -34 427589
rect 34 427555 50 427589
rect -50 427539 50 427555
rect -50 427481 50 427497
rect -50 427447 -34 427481
rect 34 427447 50 427481
rect -50 427409 50 427447
rect -50 426371 50 426409
rect -50 426337 -34 426371
rect 34 426337 50 426371
rect -50 426321 50 426337
rect -50 426263 50 426279
rect -50 426229 -34 426263
rect 34 426229 50 426263
rect -50 426191 50 426229
rect -50 425153 50 425191
rect -50 425119 -34 425153
rect 34 425119 50 425153
rect -50 425103 50 425119
rect -50 425045 50 425061
rect -50 425011 -34 425045
rect 34 425011 50 425045
rect -50 424973 50 425011
rect -50 423935 50 423973
rect -50 423901 -34 423935
rect 34 423901 50 423935
rect -50 423885 50 423901
rect -50 423827 50 423843
rect -50 423793 -34 423827
rect 34 423793 50 423827
rect -50 423755 50 423793
rect -50 422717 50 422755
rect -50 422683 -34 422717
rect 34 422683 50 422717
rect -50 422667 50 422683
rect -50 422609 50 422625
rect -50 422575 -34 422609
rect 34 422575 50 422609
rect -50 422537 50 422575
rect -50 421499 50 421537
rect -50 421465 -34 421499
rect 34 421465 50 421499
rect -50 421449 50 421465
rect -50 421391 50 421407
rect -50 421357 -34 421391
rect 34 421357 50 421391
rect -50 421319 50 421357
rect -50 420281 50 420319
rect -50 420247 -34 420281
rect 34 420247 50 420281
rect -50 420231 50 420247
rect -50 420173 50 420189
rect -50 420139 -34 420173
rect 34 420139 50 420173
rect -50 420101 50 420139
rect -50 419063 50 419101
rect -50 419029 -34 419063
rect 34 419029 50 419063
rect -50 419013 50 419029
rect -50 418955 50 418971
rect -50 418921 -34 418955
rect 34 418921 50 418955
rect -50 418883 50 418921
rect -50 417845 50 417883
rect -50 417811 -34 417845
rect 34 417811 50 417845
rect -50 417795 50 417811
rect -50 417737 50 417753
rect -50 417703 -34 417737
rect 34 417703 50 417737
rect -50 417665 50 417703
rect -50 416627 50 416665
rect -50 416593 -34 416627
rect 34 416593 50 416627
rect -50 416577 50 416593
rect -50 416519 50 416535
rect -50 416485 -34 416519
rect 34 416485 50 416519
rect -50 416447 50 416485
rect -50 415409 50 415447
rect -50 415375 -34 415409
rect 34 415375 50 415409
rect -50 415359 50 415375
rect -50 415301 50 415317
rect -50 415267 -34 415301
rect 34 415267 50 415301
rect -50 415229 50 415267
rect -50 414191 50 414229
rect -50 414157 -34 414191
rect 34 414157 50 414191
rect -50 414141 50 414157
rect -50 414083 50 414099
rect -50 414049 -34 414083
rect 34 414049 50 414083
rect -50 414011 50 414049
rect -50 412973 50 413011
rect -50 412939 -34 412973
rect 34 412939 50 412973
rect -50 412923 50 412939
rect -50 412865 50 412881
rect -50 412831 -34 412865
rect 34 412831 50 412865
rect -50 412793 50 412831
rect -50 411755 50 411793
rect -50 411721 -34 411755
rect 34 411721 50 411755
rect -50 411705 50 411721
rect -50 411647 50 411663
rect -50 411613 -34 411647
rect 34 411613 50 411647
rect -50 411575 50 411613
rect -50 410537 50 410575
rect -50 410503 -34 410537
rect 34 410503 50 410537
rect -50 410487 50 410503
rect -50 410429 50 410445
rect -50 410395 -34 410429
rect 34 410395 50 410429
rect -50 410357 50 410395
rect -50 409319 50 409357
rect -50 409285 -34 409319
rect 34 409285 50 409319
rect -50 409269 50 409285
rect -50 409211 50 409227
rect -50 409177 -34 409211
rect 34 409177 50 409211
rect -50 409139 50 409177
rect -50 408101 50 408139
rect -50 408067 -34 408101
rect 34 408067 50 408101
rect -50 408051 50 408067
rect -50 407993 50 408009
rect -50 407959 -34 407993
rect 34 407959 50 407993
rect -50 407921 50 407959
rect -50 406883 50 406921
rect -50 406849 -34 406883
rect 34 406849 50 406883
rect -50 406833 50 406849
rect -50 406775 50 406791
rect -50 406741 -34 406775
rect 34 406741 50 406775
rect -50 406703 50 406741
rect -50 405665 50 405703
rect -50 405631 -34 405665
rect 34 405631 50 405665
rect -50 405615 50 405631
rect -50 405557 50 405573
rect -50 405523 -34 405557
rect 34 405523 50 405557
rect -50 405485 50 405523
rect -50 404447 50 404485
rect -50 404413 -34 404447
rect 34 404413 50 404447
rect -50 404397 50 404413
rect -50 404339 50 404355
rect -50 404305 -34 404339
rect 34 404305 50 404339
rect -50 404267 50 404305
rect -50 403229 50 403267
rect -50 403195 -34 403229
rect 34 403195 50 403229
rect -50 403179 50 403195
rect -50 403121 50 403137
rect -50 403087 -34 403121
rect 34 403087 50 403121
rect -50 403049 50 403087
rect -50 402011 50 402049
rect -50 401977 -34 402011
rect 34 401977 50 402011
rect -50 401961 50 401977
rect -50 401903 50 401919
rect -50 401869 -34 401903
rect 34 401869 50 401903
rect -50 401831 50 401869
rect -50 400793 50 400831
rect -50 400759 -34 400793
rect 34 400759 50 400793
rect -50 400743 50 400759
rect -50 400685 50 400701
rect -50 400651 -34 400685
rect 34 400651 50 400685
rect -50 400613 50 400651
rect -50 399575 50 399613
rect -50 399541 -34 399575
rect 34 399541 50 399575
rect -50 399525 50 399541
rect -50 399467 50 399483
rect -50 399433 -34 399467
rect 34 399433 50 399467
rect -50 399395 50 399433
rect -50 398357 50 398395
rect -50 398323 -34 398357
rect 34 398323 50 398357
rect -50 398307 50 398323
rect -50 398249 50 398265
rect -50 398215 -34 398249
rect 34 398215 50 398249
rect -50 398177 50 398215
rect -50 397139 50 397177
rect -50 397105 -34 397139
rect 34 397105 50 397139
rect -50 397089 50 397105
rect -50 397031 50 397047
rect -50 396997 -34 397031
rect 34 396997 50 397031
rect -50 396959 50 396997
rect -50 395921 50 395959
rect -50 395887 -34 395921
rect 34 395887 50 395921
rect -50 395871 50 395887
rect -50 395813 50 395829
rect -50 395779 -34 395813
rect 34 395779 50 395813
rect -50 395741 50 395779
rect -50 394703 50 394741
rect -50 394669 -34 394703
rect 34 394669 50 394703
rect -50 394653 50 394669
rect -50 394595 50 394611
rect -50 394561 -34 394595
rect 34 394561 50 394595
rect -50 394523 50 394561
rect -50 393485 50 393523
rect -50 393451 -34 393485
rect 34 393451 50 393485
rect -50 393435 50 393451
rect -50 393377 50 393393
rect -50 393343 -34 393377
rect 34 393343 50 393377
rect -50 393305 50 393343
rect -50 392267 50 392305
rect -50 392233 -34 392267
rect 34 392233 50 392267
rect -50 392217 50 392233
rect -50 392159 50 392175
rect -50 392125 -34 392159
rect 34 392125 50 392159
rect -50 392087 50 392125
rect -50 391049 50 391087
rect -50 391015 -34 391049
rect 34 391015 50 391049
rect -50 390999 50 391015
rect -50 390941 50 390957
rect -50 390907 -34 390941
rect 34 390907 50 390941
rect -50 390869 50 390907
rect -50 389831 50 389869
rect -50 389797 -34 389831
rect 34 389797 50 389831
rect -50 389781 50 389797
rect -50 389723 50 389739
rect -50 389689 -34 389723
rect 34 389689 50 389723
rect -50 389651 50 389689
rect -50 388613 50 388651
rect -50 388579 -34 388613
rect 34 388579 50 388613
rect -50 388563 50 388579
rect -50 388505 50 388521
rect -50 388471 -34 388505
rect 34 388471 50 388505
rect -50 388433 50 388471
rect -50 387395 50 387433
rect -50 387361 -34 387395
rect 34 387361 50 387395
rect -50 387345 50 387361
rect -50 387287 50 387303
rect -50 387253 -34 387287
rect 34 387253 50 387287
rect -50 387215 50 387253
rect -50 386177 50 386215
rect -50 386143 -34 386177
rect 34 386143 50 386177
rect -50 386127 50 386143
rect -50 386069 50 386085
rect -50 386035 -34 386069
rect 34 386035 50 386069
rect -50 385997 50 386035
rect -50 384959 50 384997
rect -50 384925 -34 384959
rect 34 384925 50 384959
rect -50 384909 50 384925
rect -50 384851 50 384867
rect -50 384817 -34 384851
rect 34 384817 50 384851
rect -50 384779 50 384817
rect -50 383741 50 383779
rect -50 383707 -34 383741
rect 34 383707 50 383741
rect -50 383691 50 383707
rect -50 383633 50 383649
rect -50 383599 -34 383633
rect 34 383599 50 383633
rect -50 383561 50 383599
rect -50 382523 50 382561
rect -50 382489 -34 382523
rect 34 382489 50 382523
rect -50 382473 50 382489
rect -50 382415 50 382431
rect -50 382381 -34 382415
rect 34 382381 50 382415
rect -50 382343 50 382381
rect -50 381305 50 381343
rect -50 381271 -34 381305
rect 34 381271 50 381305
rect -50 381255 50 381271
rect -50 381197 50 381213
rect -50 381163 -34 381197
rect 34 381163 50 381197
rect -50 381125 50 381163
rect -50 380087 50 380125
rect -50 380053 -34 380087
rect 34 380053 50 380087
rect -50 380037 50 380053
rect -50 379979 50 379995
rect -50 379945 -34 379979
rect 34 379945 50 379979
rect -50 379907 50 379945
rect -50 378869 50 378907
rect -50 378835 -34 378869
rect 34 378835 50 378869
rect -50 378819 50 378835
rect -50 378761 50 378777
rect -50 378727 -34 378761
rect 34 378727 50 378761
rect -50 378689 50 378727
rect -50 377651 50 377689
rect -50 377617 -34 377651
rect 34 377617 50 377651
rect -50 377601 50 377617
rect -50 377543 50 377559
rect -50 377509 -34 377543
rect 34 377509 50 377543
rect -50 377471 50 377509
rect -50 376433 50 376471
rect -50 376399 -34 376433
rect 34 376399 50 376433
rect -50 376383 50 376399
rect -50 376325 50 376341
rect -50 376291 -34 376325
rect 34 376291 50 376325
rect -50 376253 50 376291
rect -50 375215 50 375253
rect -50 375181 -34 375215
rect 34 375181 50 375215
rect -50 375165 50 375181
rect -50 375107 50 375123
rect -50 375073 -34 375107
rect 34 375073 50 375107
rect -50 375035 50 375073
rect -50 373997 50 374035
rect -50 373963 -34 373997
rect 34 373963 50 373997
rect -50 373947 50 373963
rect -50 373889 50 373905
rect -50 373855 -34 373889
rect 34 373855 50 373889
rect -50 373817 50 373855
rect -50 372779 50 372817
rect -50 372745 -34 372779
rect 34 372745 50 372779
rect -50 372729 50 372745
rect -50 372671 50 372687
rect -50 372637 -34 372671
rect 34 372637 50 372671
rect -50 372599 50 372637
rect -50 371561 50 371599
rect -50 371527 -34 371561
rect 34 371527 50 371561
rect -50 371511 50 371527
rect -50 371453 50 371469
rect -50 371419 -34 371453
rect 34 371419 50 371453
rect -50 371381 50 371419
rect -50 370343 50 370381
rect -50 370309 -34 370343
rect 34 370309 50 370343
rect -50 370293 50 370309
rect -50 370235 50 370251
rect -50 370201 -34 370235
rect 34 370201 50 370235
rect -50 370163 50 370201
rect -50 369125 50 369163
rect -50 369091 -34 369125
rect 34 369091 50 369125
rect -50 369075 50 369091
rect -50 369017 50 369033
rect -50 368983 -34 369017
rect 34 368983 50 369017
rect -50 368945 50 368983
rect -50 367907 50 367945
rect -50 367873 -34 367907
rect 34 367873 50 367907
rect -50 367857 50 367873
rect -50 367799 50 367815
rect -50 367765 -34 367799
rect 34 367765 50 367799
rect -50 367727 50 367765
rect -50 366689 50 366727
rect -50 366655 -34 366689
rect 34 366655 50 366689
rect -50 366639 50 366655
rect -50 366581 50 366597
rect -50 366547 -34 366581
rect 34 366547 50 366581
rect -50 366509 50 366547
rect -50 365471 50 365509
rect -50 365437 -34 365471
rect 34 365437 50 365471
rect -50 365421 50 365437
rect -50 365363 50 365379
rect -50 365329 -34 365363
rect 34 365329 50 365363
rect -50 365291 50 365329
rect -50 364253 50 364291
rect -50 364219 -34 364253
rect 34 364219 50 364253
rect -50 364203 50 364219
rect -50 364145 50 364161
rect -50 364111 -34 364145
rect 34 364111 50 364145
rect -50 364073 50 364111
rect -50 363035 50 363073
rect -50 363001 -34 363035
rect 34 363001 50 363035
rect -50 362985 50 363001
rect -50 362927 50 362943
rect -50 362893 -34 362927
rect 34 362893 50 362927
rect -50 362855 50 362893
rect -50 361817 50 361855
rect -50 361783 -34 361817
rect 34 361783 50 361817
rect -50 361767 50 361783
rect -50 361709 50 361725
rect -50 361675 -34 361709
rect 34 361675 50 361709
rect -50 361637 50 361675
rect -50 360599 50 360637
rect -50 360565 -34 360599
rect 34 360565 50 360599
rect -50 360549 50 360565
rect -50 360491 50 360507
rect -50 360457 -34 360491
rect 34 360457 50 360491
rect -50 360419 50 360457
rect -50 359381 50 359419
rect -50 359347 -34 359381
rect 34 359347 50 359381
rect -50 359331 50 359347
rect -50 359273 50 359289
rect -50 359239 -34 359273
rect 34 359239 50 359273
rect -50 359201 50 359239
rect -50 358163 50 358201
rect -50 358129 -34 358163
rect 34 358129 50 358163
rect -50 358113 50 358129
rect -50 358055 50 358071
rect -50 358021 -34 358055
rect 34 358021 50 358055
rect -50 357983 50 358021
rect -50 356945 50 356983
rect -50 356911 -34 356945
rect 34 356911 50 356945
rect -50 356895 50 356911
rect -50 356837 50 356853
rect -50 356803 -34 356837
rect 34 356803 50 356837
rect -50 356765 50 356803
rect -50 355727 50 355765
rect -50 355693 -34 355727
rect 34 355693 50 355727
rect -50 355677 50 355693
rect -50 355619 50 355635
rect -50 355585 -34 355619
rect 34 355585 50 355619
rect -50 355547 50 355585
rect -50 354509 50 354547
rect -50 354475 -34 354509
rect 34 354475 50 354509
rect -50 354459 50 354475
rect -50 354401 50 354417
rect -50 354367 -34 354401
rect 34 354367 50 354401
rect -50 354329 50 354367
rect -50 353291 50 353329
rect -50 353257 -34 353291
rect 34 353257 50 353291
rect -50 353241 50 353257
rect -50 353183 50 353199
rect -50 353149 -34 353183
rect 34 353149 50 353183
rect -50 353111 50 353149
rect -50 352073 50 352111
rect -50 352039 -34 352073
rect 34 352039 50 352073
rect -50 352023 50 352039
rect -50 351965 50 351981
rect -50 351931 -34 351965
rect 34 351931 50 351965
rect -50 351893 50 351931
rect -50 350855 50 350893
rect -50 350821 -34 350855
rect 34 350821 50 350855
rect -50 350805 50 350821
rect -50 350747 50 350763
rect -50 350713 -34 350747
rect 34 350713 50 350747
rect -50 350675 50 350713
rect -50 349637 50 349675
rect -50 349603 -34 349637
rect 34 349603 50 349637
rect -50 349587 50 349603
rect -50 349529 50 349545
rect -50 349495 -34 349529
rect 34 349495 50 349529
rect -50 349457 50 349495
rect -50 348419 50 348457
rect -50 348385 -34 348419
rect 34 348385 50 348419
rect -50 348369 50 348385
rect -50 348311 50 348327
rect -50 348277 -34 348311
rect 34 348277 50 348311
rect -50 348239 50 348277
rect -50 347201 50 347239
rect -50 347167 -34 347201
rect 34 347167 50 347201
rect -50 347151 50 347167
rect -50 347093 50 347109
rect -50 347059 -34 347093
rect 34 347059 50 347093
rect -50 347021 50 347059
rect -50 345983 50 346021
rect -50 345949 -34 345983
rect 34 345949 50 345983
rect -50 345933 50 345949
rect -50 345875 50 345891
rect -50 345841 -34 345875
rect 34 345841 50 345875
rect -50 345803 50 345841
rect -50 344765 50 344803
rect -50 344731 -34 344765
rect 34 344731 50 344765
rect -50 344715 50 344731
rect -50 344657 50 344673
rect -50 344623 -34 344657
rect 34 344623 50 344657
rect -50 344585 50 344623
rect -50 343547 50 343585
rect -50 343513 -34 343547
rect 34 343513 50 343547
rect -50 343497 50 343513
rect -50 343439 50 343455
rect -50 343405 -34 343439
rect 34 343405 50 343439
rect -50 343367 50 343405
rect -50 342329 50 342367
rect -50 342295 -34 342329
rect 34 342295 50 342329
rect -50 342279 50 342295
rect -50 342221 50 342237
rect -50 342187 -34 342221
rect 34 342187 50 342221
rect -50 342149 50 342187
rect -50 341111 50 341149
rect -50 341077 -34 341111
rect 34 341077 50 341111
rect -50 341061 50 341077
rect -50 341003 50 341019
rect -50 340969 -34 341003
rect 34 340969 50 341003
rect -50 340931 50 340969
rect -50 339893 50 339931
rect -50 339859 -34 339893
rect 34 339859 50 339893
rect -50 339843 50 339859
rect -50 339785 50 339801
rect -50 339751 -34 339785
rect 34 339751 50 339785
rect -50 339713 50 339751
rect -50 338675 50 338713
rect -50 338641 -34 338675
rect 34 338641 50 338675
rect -50 338625 50 338641
rect -50 338567 50 338583
rect -50 338533 -34 338567
rect 34 338533 50 338567
rect -50 338495 50 338533
rect -50 337457 50 337495
rect -50 337423 -34 337457
rect 34 337423 50 337457
rect -50 337407 50 337423
rect -50 337349 50 337365
rect -50 337315 -34 337349
rect 34 337315 50 337349
rect -50 337277 50 337315
rect -50 336239 50 336277
rect -50 336205 -34 336239
rect 34 336205 50 336239
rect -50 336189 50 336205
rect -50 336131 50 336147
rect -50 336097 -34 336131
rect 34 336097 50 336131
rect -50 336059 50 336097
rect -50 335021 50 335059
rect -50 334987 -34 335021
rect 34 334987 50 335021
rect -50 334971 50 334987
rect -50 334913 50 334929
rect -50 334879 -34 334913
rect 34 334879 50 334913
rect -50 334841 50 334879
rect -50 333803 50 333841
rect -50 333769 -34 333803
rect 34 333769 50 333803
rect -50 333753 50 333769
rect -50 333695 50 333711
rect -50 333661 -34 333695
rect 34 333661 50 333695
rect -50 333623 50 333661
rect -50 332585 50 332623
rect -50 332551 -34 332585
rect 34 332551 50 332585
rect -50 332535 50 332551
rect -50 332477 50 332493
rect -50 332443 -34 332477
rect 34 332443 50 332477
rect -50 332405 50 332443
rect -50 331367 50 331405
rect -50 331333 -34 331367
rect 34 331333 50 331367
rect -50 331317 50 331333
rect -50 331259 50 331275
rect -50 331225 -34 331259
rect 34 331225 50 331259
rect -50 331187 50 331225
rect -50 330149 50 330187
rect -50 330115 -34 330149
rect 34 330115 50 330149
rect -50 330099 50 330115
rect -50 330041 50 330057
rect -50 330007 -34 330041
rect 34 330007 50 330041
rect -50 329969 50 330007
rect -50 328931 50 328969
rect -50 328897 -34 328931
rect 34 328897 50 328931
rect -50 328881 50 328897
rect -50 328823 50 328839
rect -50 328789 -34 328823
rect 34 328789 50 328823
rect -50 328751 50 328789
rect -50 327713 50 327751
rect -50 327679 -34 327713
rect 34 327679 50 327713
rect -50 327663 50 327679
rect -50 327605 50 327621
rect -50 327571 -34 327605
rect 34 327571 50 327605
rect -50 327533 50 327571
rect -50 326495 50 326533
rect -50 326461 -34 326495
rect 34 326461 50 326495
rect -50 326445 50 326461
rect -50 326387 50 326403
rect -50 326353 -34 326387
rect 34 326353 50 326387
rect -50 326315 50 326353
rect -50 325277 50 325315
rect -50 325243 -34 325277
rect 34 325243 50 325277
rect -50 325227 50 325243
rect -50 325169 50 325185
rect -50 325135 -34 325169
rect 34 325135 50 325169
rect -50 325097 50 325135
rect -50 324059 50 324097
rect -50 324025 -34 324059
rect 34 324025 50 324059
rect -50 324009 50 324025
rect -50 323951 50 323967
rect -50 323917 -34 323951
rect 34 323917 50 323951
rect -50 323879 50 323917
rect -50 322841 50 322879
rect -50 322807 -34 322841
rect 34 322807 50 322841
rect -50 322791 50 322807
rect -50 322733 50 322749
rect -50 322699 -34 322733
rect 34 322699 50 322733
rect -50 322661 50 322699
rect -50 321623 50 321661
rect -50 321589 -34 321623
rect 34 321589 50 321623
rect -50 321573 50 321589
rect -50 321515 50 321531
rect -50 321481 -34 321515
rect 34 321481 50 321515
rect -50 321443 50 321481
rect -50 320405 50 320443
rect -50 320371 -34 320405
rect 34 320371 50 320405
rect -50 320355 50 320371
rect -50 320297 50 320313
rect -50 320263 -34 320297
rect 34 320263 50 320297
rect -50 320225 50 320263
rect -50 319187 50 319225
rect -50 319153 -34 319187
rect 34 319153 50 319187
rect -50 319137 50 319153
rect -50 319079 50 319095
rect -50 319045 -34 319079
rect 34 319045 50 319079
rect -50 319007 50 319045
rect -50 317969 50 318007
rect -50 317935 -34 317969
rect 34 317935 50 317969
rect -50 317919 50 317935
rect -50 317861 50 317877
rect -50 317827 -34 317861
rect 34 317827 50 317861
rect -50 317789 50 317827
rect -50 316751 50 316789
rect -50 316717 -34 316751
rect 34 316717 50 316751
rect -50 316701 50 316717
rect -50 316643 50 316659
rect -50 316609 -34 316643
rect 34 316609 50 316643
rect -50 316571 50 316609
rect -50 315533 50 315571
rect -50 315499 -34 315533
rect 34 315499 50 315533
rect -50 315483 50 315499
rect -50 315425 50 315441
rect -50 315391 -34 315425
rect 34 315391 50 315425
rect -50 315353 50 315391
rect -50 314315 50 314353
rect -50 314281 -34 314315
rect 34 314281 50 314315
rect -50 314265 50 314281
rect -50 314207 50 314223
rect -50 314173 -34 314207
rect 34 314173 50 314207
rect -50 314135 50 314173
rect -50 313097 50 313135
rect -50 313063 -34 313097
rect 34 313063 50 313097
rect -50 313047 50 313063
rect -50 312989 50 313005
rect -50 312955 -34 312989
rect 34 312955 50 312989
rect -50 312917 50 312955
rect -50 311879 50 311917
rect -50 311845 -34 311879
rect 34 311845 50 311879
rect -50 311829 50 311845
rect -50 311771 50 311787
rect -50 311737 -34 311771
rect 34 311737 50 311771
rect -50 311699 50 311737
rect -50 310661 50 310699
rect -50 310627 -34 310661
rect 34 310627 50 310661
rect -50 310611 50 310627
rect -50 310553 50 310569
rect -50 310519 -34 310553
rect 34 310519 50 310553
rect -50 310481 50 310519
rect -50 309443 50 309481
rect -50 309409 -34 309443
rect 34 309409 50 309443
rect -50 309393 50 309409
rect -50 309335 50 309351
rect -50 309301 -34 309335
rect 34 309301 50 309335
rect -50 309263 50 309301
rect -50 308225 50 308263
rect -50 308191 -34 308225
rect 34 308191 50 308225
rect -50 308175 50 308191
rect -50 308117 50 308133
rect -50 308083 -34 308117
rect 34 308083 50 308117
rect -50 308045 50 308083
rect -50 307007 50 307045
rect -50 306973 -34 307007
rect 34 306973 50 307007
rect -50 306957 50 306973
rect -50 306899 50 306915
rect -50 306865 -34 306899
rect 34 306865 50 306899
rect -50 306827 50 306865
rect -50 305789 50 305827
rect -50 305755 -34 305789
rect 34 305755 50 305789
rect -50 305739 50 305755
rect -50 305681 50 305697
rect -50 305647 -34 305681
rect 34 305647 50 305681
rect -50 305609 50 305647
rect -50 304571 50 304609
rect -50 304537 -34 304571
rect 34 304537 50 304571
rect -50 304521 50 304537
rect -50 304463 50 304479
rect -50 304429 -34 304463
rect 34 304429 50 304463
rect -50 304391 50 304429
rect -50 303353 50 303391
rect -50 303319 -34 303353
rect 34 303319 50 303353
rect -50 303303 50 303319
rect -50 303245 50 303261
rect -50 303211 -34 303245
rect 34 303211 50 303245
rect -50 303173 50 303211
rect -50 302135 50 302173
rect -50 302101 -34 302135
rect 34 302101 50 302135
rect -50 302085 50 302101
rect -50 302027 50 302043
rect -50 301993 -34 302027
rect 34 301993 50 302027
rect -50 301955 50 301993
rect -50 300917 50 300955
rect -50 300883 -34 300917
rect 34 300883 50 300917
rect -50 300867 50 300883
rect -50 300809 50 300825
rect -50 300775 -34 300809
rect 34 300775 50 300809
rect -50 300737 50 300775
rect -50 299699 50 299737
rect -50 299665 -34 299699
rect 34 299665 50 299699
rect -50 299649 50 299665
rect -50 299591 50 299607
rect -50 299557 -34 299591
rect 34 299557 50 299591
rect -50 299519 50 299557
rect -50 298481 50 298519
rect -50 298447 -34 298481
rect 34 298447 50 298481
rect -50 298431 50 298447
rect -50 298373 50 298389
rect -50 298339 -34 298373
rect 34 298339 50 298373
rect -50 298301 50 298339
rect -50 297263 50 297301
rect -50 297229 -34 297263
rect 34 297229 50 297263
rect -50 297213 50 297229
rect -50 297155 50 297171
rect -50 297121 -34 297155
rect 34 297121 50 297155
rect -50 297083 50 297121
rect -50 296045 50 296083
rect -50 296011 -34 296045
rect 34 296011 50 296045
rect -50 295995 50 296011
rect -50 295937 50 295953
rect -50 295903 -34 295937
rect 34 295903 50 295937
rect -50 295865 50 295903
rect -50 294827 50 294865
rect -50 294793 -34 294827
rect 34 294793 50 294827
rect -50 294777 50 294793
rect -50 294719 50 294735
rect -50 294685 -34 294719
rect 34 294685 50 294719
rect -50 294647 50 294685
rect -50 293609 50 293647
rect -50 293575 -34 293609
rect 34 293575 50 293609
rect -50 293559 50 293575
rect -50 293501 50 293517
rect -50 293467 -34 293501
rect 34 293467 50 293501
rect -50 293429 50 293467
rect -50 292391 50 292429
rect -50 292357 -34 292391
rect 34 292357 50 292391
rect -50 292341 50 292357
rect -50 292283 50 292299
rect -50 292249 -34 292283
rect 34 292249 50 292283
rect -50 292211 50 292249
rect -50 291173 50 291211
rect -50 291139 -34 291173
rect 34 291139 50 291173
rect -50 291123 50 291139
rect -50 291065 50 291081
rect -50 291031 -34 291065
rect 34 291031 50 291065
rect -50 290993 50 291031
rect -50 289955 50 289993
rect -50 289921 -34 289955
rect 34 289921 50 289955
rect -50 289905 50 289921
rect -50 289847 50 289863
rect -50 289813 -34 289847
rect 34 289813 50 289847
rect -50 289775 50 289813
rect -50 288737 50 288775
rect -50 288703 -34 288737
rect 34 288703 50 288737
rect -50 288687 50 288703
rect -50 288629 50 288645
rect -50 288595 -34 288629
rect 34 288595 50 288629
rect -50 288557 50 288595
rect -50 287519 50 287557
rect -50 287485 -34 287519
rect 34 287485 50 287519
rect -50 287469 50 287485
rect -50 287411 50 287427
rect -50 287377 -34 287411
rect 34 287377 50 287411
rect -50 287339 50 287377
rect -50 286301 50 286339
rect -50 286267 -34 286301
rect 34 286267 50 286301
rect -50 286251 50 286267
rect -50 286193 50 286209
rect -50 286159 -34 286193
rect 34 286159 50 286193
rect -50 286121 50 286159
rect -50 285083 50 285121
rect -50 285049 -34 285083
rect 34 285049 50 285083
rect -50 285033 50 285049
rect -50 284975 50 284991
rect -50 284941 -34 284975
rect 34 284941 50 284975
rect -50 284903 50 284941
rect -50 283865 50 283903
rect -50 283831 -34 283865
rect 34 283831 50 283865
rect -50 283815 50 283831
rect -50 283757 50 283773
rect -50 283723 -34 283757
rect 34 283723 50 283757
rect -50 283685 50 283723
rect -50 282647 50 282685
rect -50 282613 -34 282647
rect 34 282613 50 282647
rect -50 282597 50 282613
rect -50 282539 50 282555
rect -50 282505 -34 282539
rect 34 282505 50 282539
rect -50 282467 50 282505
rect -50 281429 50 281467
rect -50 281395 -34 281429
rect 34 281395 50 281429
rect -50 281379 50 281395
rect -50 281321 50 281337
rect -50 281287 -34 281321
rect 34 281287 50 281321
rect -50 281249 50 281287
rect -50 280211 50 280249
rect -50 280177 -34 280211
rect 34 280177 50 280211
rect -50 280161 50 280177
rect -50 280103 50 280119
rect -50 280069 -34 280103
rect 34 280069 50 280103
rect -50 280031 50 280069
rect -50 278993 50 279031
rect -50 278959 -34 278993
rect 34 278959 50 278993
rect -50 278943 50 278959
rect -50 278885 50 278901
rect -50 278851 -34 278885
rect 34 278851 50 278885
rect -50 278813 50 278851
rect -50 277775 50 277813
rect -50 277741 -34 277775
rect 34 277741 50 277775
rect -50 277725 50 277741
rect -50 277667 50 277683
rect -50 277633 -34 277667
rect 34 277633 50 277667
rect -50 277595 50 277633
rect -50 276557 50 276595
rect -50 276523 -34 276557
rect 34 276523 50 276557
rect -50 276507 50 276523
rect -50 276449 50 276465
rect -50 276415 -34 276449
rect 34 276415 50 276449
rect -50 276377 50 276415
rect -50 275339 50 275377
rect -50 275305 -34 275339
rect 34 275305 50 275339
rect -50 275289 50 275305
rect -50 275231 50 275247
rect -50 275197 -34 275231
rect 34 275197 50 275231
rect -50 275159 50 275197
rect -50 274121 50 274159
rect -50 274087 -34 274121
rect 34 274087 50 274121
rect -50 274071 50 274087
rect -50 274013 50 274029
rect -50 273979 -34 274013
rect 34 273979 50 274013
rect -50 273941 50 273979
rect -50 272903 50 272941
rect -50 272869 -34 272903
rect 34 272869 50 272903
rect -50 272853 50 272869
rect -50 272795 50 272811
rect -50 272761 -34 272795
rect 34 272761 50 272795
rect -50 272723 50 272761
rect -50 271685 50 271723
rect -50 271651 -34 271685
rect 34 271651 50 271685
rect -50 271635 50 271651
rect -50 271577 50 271593
rect -50 271543 -34 271577
rect 34 271543 50 271577
rect -50 271505 50 271543
rect -50 270467 50 270505
rect -50 270433 -34 270467
rect 34 270433 50 270467
rect -50 270417 50 270433
rect -50 270359 50 270375
rect -50 270325 -34 270359
rect 34 270325 50 270359
rect -50 270287 50 270325
rect -50 269249 50 269287
rect -50 269215 -34 269249
rect 34 269215 50 269249
rect -50 269199 50 269215
rect -50 269141 50 269157
rect -50 269107 -34 269141
rect 34 269107 50 269141
rect -50 269069 50 269107
rect -50 268031 50 268069
rect -50 267997 -34 268031
rect 34 267997 50 268031
rect -50 267981 50 267997
rect -50 267923 50 267939
rect -50 267889 -34 267923
rect 34 267889 50 267923
rect -50 267851 50 267889
rect -50 266813 50 266851
rect -50 266779 -34 266813
rect 34 266779 50 266813
rect -50 266763 50 266779
rect -50 266705 50 266721
rect -50 266671 -34 266705
rect 34 266671 50 266705
rect -50 266633 50 266671
rect -50 265595 50 265633
rect -50 265561 -34 265595
rect 34 265561 50 265595
rect -50 265545 50 265561
rect -50 265487 50 265503
rect -50 265453 -34 265487
rect 34 265453 50 265487
rect -50 265415 50 265453
rect -50 264377 50 264415
rect -50 264343 -34 264377
rect 34 264343 50 264377
rect -50 264327 50 264343
rect -50 264269 50 264285
rect -50 264235 -34 264269
rect 34 264235 50 264269
rect -50 264197 50 264235
rect -50 263159 50 263197
rect -50 263125 -34 263159
rect 34 263125 50 263159
rect -50 263109 50 263125
rect -50 263051 50 263067
rect -50 263017 -34 263051
rect 34 263017 50 263051
rect -50 262979 50 263017
rect -50 261941 50 261979
rect -50 261907 -34 261941
rect 34 261907 50 261941
rect -50 261891 50 261907
rect -50 261833 50 261849
rect -50 261799 -34 261833
rect 34 261799 50 261833
rect -50 261761 50 261799
rect -50 260723 50 260761
rect -50 260689 -34 260723
rect 34 260689 50 260723
rect -50 260673 50 260689
rect -50 260615 50 260631
rect -50 260581 -34 260615
rect 34 260581 50 260615
rect -50 260543 50 260581
rect -50 259505 50 259543
rect -50 259471 -34 259505
rect 34 259471 50 259505
rect -50 259455 50 259471
rect -50 259397 50 259413
rect -50 259363 -34 259397
rect 34 259363 50 259397
rect -50 259325 50 259363
rect -50 258287 50 258325
rect -50 258253 -34 258287
rect 34 258253 50 258287
rect -50 258237 50 258253
rect -50 258179 50 258195
rect -50 258145 -34 258179
rect 34 258145 50 258179
rect -50 258107 50 258145
rect -50 257069 50 257107
rect -50 257035 -34 257069
rect 34 257035 50 257069
rect -50 257019 50 257035
rect -50 256961 50 256977
rect -50 256927 -34 256961
rect 34 256927 50 256961
rect -50 256889 50 256927
rect -50 255851 50 255889
rect -50 255817 -34 255851
rect 34 255817 50 255851
rect -50 255801 50 255817
rect -50 255743 50 255759
rect -50 255709 -34 255743
rect 34 255709 50 255743
rect -50 255671 50 255709
rect -50 254633 50 254671
rect -50 254599 -34 254633
rect 34 254599 50 254633
rect -50 254583 50 254599
rect -50 254525 50 254541
rect -50 254491 -34 254525
rect 34 254491 50 254525
rect -50 254453 50 254491
rect -50 253415 50 253453
rect -50 253381 -34 253415
rect 34 253381 50 253415
rect -50 253365 50 253381
rect -50 253307 50 253323
rect -50 253273 -34 253307
rect 34 253273 50 253307
rect -50 253235 50 253273
rect -50 252197 50 252235
rect -50 252163 -34 252197
rect 34 252163 50 252197
rect -50 252147 50 252163
rect -50 252089 50 252105
rect -50 252055 -34 252089
rect 34 252055 50 252089
rect -50 252017 50 252055
rect -50 250979 50 251017
rect -50 250945 -34 250979
rect 34 250945 50 250979
rect -50 250929 50 250945
rect -50 250871 50 250887
rect -50 250837 -34 250871
rect 34 250837 50 250871
rect -50 250799 50 250837
rect -50 249761 50 249799
rect -50 249727 -34 249761
rect 34 249727 50 249761
rect -50 249711 50 249727
rect -50 249653 50 249669
rect -50 249619 -34 249653
rect 34 249619 50 249653
rect -50 249581 50 249619
rect -50 248543 50 248581
rect -50 248509 -34 248543
rect 34 248509 50 248543
rect -50 248493 50 248509
rect -50 248435 50 248451
rect -50 248401 -34 248435
rect 34 248401 50 248435
rect -50 248363 50 248401
rect -50 247325 50 247363
rect -50 247291 -34 247325
rect 34 247291 50 247325
rect -50 247275 50 247291
rect -50 247217 50 247233
rect -50 247183 -34 247217
rect 34 247183 50 247217
rect -50 247145 50 247183
rect -50 246107 50 246145
rect -50 246073 -34 246107
rect 34 246073 50 246107
rect -50 246057 50 246073
rect -50 245999 50 246015
rect -50 245965 -34 245999
rect 34 245965 50 245999
rect -50 245927 50 245965
rect -50 244889 50 244927
rect -50 244855 -34 244889
rect 34 244855 50 244889
rect -50 244839 50 244855
rect -50 244781 50 244797
rect -50 244747 -34 244781
rect 34 244747 50 244781
rect -50 244709 50 244747
rect -50 243671 50 243709
rect -50 243637 -34 243671
rect 34 243637 50 243671
rect -50 243621 50 243637
rect -50 243563 50 243579
rect -50 243529 -34 243563
rect 34 243529 50 243563
rect -50 243491 50 243529
rect -50 242453 50 242491
rect -50 242419 -34 242453
rect 34 242419 50 242453
rect -50 242403 50 242419
rect -50 242345 50 242361
rect -50 242311 -34 242345
rect 34 242311 50 242345
rect -50 242273 50 242311
rect -50 241235 50 241273
rect -50 241201 -34 241235
rect 34 241201 50 241235
rect -50 241185 50 241201
rect -50 241127 50 241143
rect -50 241093 -34 241127
rect 34 241093 50 241127
rect -50 241055 50 241093
rect -50 240017 50 240055
rect -50 239983 -34 240017
rect 34 239983 50 240017
rect -50 239967 50 239983
rect -50 239909 50 239925
rect -50 239875 -34 239909
rect 34 239875 50 239909
rect -50 239837 50 239875
rect -50 238799 50 238837
rect -50 238765 -34 238799
rect 34 238765 50 238799
rect -50 238749 50 238765
rect -50 238691 50 238707
rect -50 238657 -34 238691
rect 34 238657 50 238691
rect -50 238619 50 238657
rect -50 237581 50 237619
rect -50 237547 -34 237581
rect 34 237547 50 237581
rect -50 237531 50 237547
rect -50 237473 50 237489
rect -50 237439 -34 237473
rect 34 237439 50 237473
rect -50 237401 50 237439
rect -50 236363 50 236401
rect -50 236329 -34 236363
rect 34 236329 50 236363
rect -50 236313 50 236329
rect -50 236255 50 236271
rect -50 236221 -34 236255
rect 34 236221 50 236255
rect -50 236183 50 236221
rect -50 235145 50 235183
rect -50 235111 -34 235145
rect 34 235111 50 235145
rect -50 235095 50 235111
rect -50 235037 50 235053
rect -50 235003 -34 235037
rect 34 235003 50 235037
rect -50 234965 50 235003
rect -50 233927 50 233965
rect -50 233893 -34 233927
rect 34 233893 50 233927
rect -50 233877 50 233893
rect -50 233819 50 233835
rect -50 233785 -34 233819
rect 34 233785 50 233819
rect -50 233747 50 233785
rect -50 232709 50 232747
rect -50 232675 -34 232709
rect 34 232675 50 232709
rect -50 232659 50 232675
rect -50 232601 50 232617
rect -50 232567 -34 232601
rect 34 232567 50 232601
rect -50 232529 50 232567
rect -50 231491 50 231529
rect -50 231457 -34 231491
rect 34 231457 50 231491
rect -50 231441 50 231457
rect -50 231383 50 231399
rect -50 231349 -34 231383
rect 34 231349 50 231383
rect -50 231311 50 231349
rect -50 230273 50 230311
rect -50 230239 -34 230273
rect 34 230239 50 230273
rect -50 230223 50 230239
rect -50 230165 50 230181
rect -50 230131 -34 230165
rect 34 230131 50 230165
rect -50 230093 50 230131
rect -50 229055 50 229093
rect -50 229021 -34 229055
rect 34 229021 50 229055
rect -50 229005 50 229021
rect -50 228947 50 228963
rect -50 228913 -34 228947
rect 34 228913 50 228947
rect -50 228875 50 228913
rect -50 227837 50 227875
rect -50 227803 -34 227837
rect 34 227803 50 227837
rect -50 227787 50 227803
rect -50 227729 50 227745
rect -50 227695 -34 227729
rect 34 227695 50 227729
rect -50 227657 50 227695
rect -50 226619 50 226657
rect -50 226585 -34 226619
rect 34 226585 50 226619
rect -50 226569 50 226585
rect -50 226511 50 226527
rect -50 226477 -34 226511
rect 34 226477 50 226511
rect -50 226439 50 226477
rect -50 225401 50 225439
rect -50 225367 -34 225401
rect 34 225367 50 225401
rect -50 225351 50 225367
rect -50 225293 50 225309
rect -50 225259 -34 225293
rect 34 225259 50 225293
rect -50 225221 50 225259
rect -50 224183 50 224221
rect -50 224149 -34 224183
rect 34 224149 50 224183
rect -50 224133 50 224149
rect -50 224075 50 224091
rect -50 224041 -34 224075
rect 34 224041 50 224075
rect -50 224003 50 224041
rect -50 222965 50 223003
rect -50 222931 -34 222965
rect 34 222931 50 222965
rect -50 222915 50 222931
rect -50 222857 50 222873
rect -50 222823 -34 222857
rect 34 222823 50 222857
rect -50 222785 50 222823
rect -50 221747 50 221785
rect -50 221713 -34 221747
rect 34 221713 50 221747
rect -50 221697 50 221713
rect -50 221639 50 221655
rect -50 221605 -34 221639
rect 34 221605 50 221639
rect -50 221567 50 221605
rect -50 220529 50 220567
rect -50 220495 -34 220529
rect 34 220495 50 220529
rect -50 220479 50 220495
rect -50 220421 50 220437
rect -50 220387 -34 220421
rect 34 220387 50 220421
rect -50 220349 50 220387
rect -50 219311 50 219349
rect -50 219277 -34 219311
rect 34 219277 50 219311
rect -50 219261 50 219277
rect -50 219203 50 219219
rect -50 219169 -34 219203
rect 34 219169 50 219203
rect -50 219131 50 219169
rect -50 218093 50 218131
rect -50 218059 -34 218093
rect 34 218059 50 218093
rect -50 218043 50 218059
rect -50 217985 50 218001
rect -50 217951 -34 217985
rect 34 217951 50 217985
rect -50 217913 50 217951
rect -50 216875 50 216913
rect -50 216841 -34 216875
rect 34 216841 50 216875
rect -50 216825 50 216841
rect -50 216767 50 216783
rect -50 216733 -34 216767
rect 34 216733 50 216767
rect -50 216695 50 216733
rect -50 215657 50 215695
rect -50 215623 -34 215657
rect 34 215623 50 215657
rect -50 215607 50 215623
rect -50 215549 50 215565
rect -50 215515 -34 215549
rect 34 215515 50 215549
rect -50 215477 50 215515
rect -50 214439 50 214477
rect -50 214405 -34 214439
rect 34 214405 50 214439
rect -50 214389 50 214405
rect -50 214331 50 214347
rect -50 214297 -34 214331
rect 34 214297 50 214331
rect -50 214259 50 214297
rect -50 213221 50 213259
rect -50 213187 -34 213221
rect 34 213187 50 213221
rect -50 213171 50 213187
rect -50 213113 50 213129
rect -50 213079 -34 213113
rect 34 213079 50 213113
rect -50 213041 50 213079
rect -50 212003 50 212041
rect -50 211969 -34 212003
rect 34 211969 50 212003
rect -50 211953 50 211969
rect -50 211895 50 211911
rect -50 211861 -34 211895
rect 34 211861 50 211895
rect -50 211823 50 211861
rect -50 210785 50 210823
rect -50 210751 -34 210785
rect 34 210751 50 210785
rect -50 210735 50 210751
rect -50 210677 50 210693
rect -50 210643 -34 210677
rect 34 210643 50 210677
rect -50 210605 50 210643
rect -50 209567 50 209605
rect -50 209533 -34 209567
rect 34 209533 50 209567
rect -50 209517 50 209533
rect -50 209459 50 209475
rect -50 209425 -34 209459
rect 34 209425 50 209459
rect -50 209387 50 209425
rect -50 208349 50 208387
rect -50 208315 -34 208349
rect 34 208315 50 208349
rect -50 208299 50 208315
rect -50 208241 50 208257
rect -50 208207 -34 208241
rect 34 208207 50 208241
rect -50 208169 50 208207
rect -50 207131 50 207169
rect -50 207097 -34 207131
rect 34 207097 50 207131
rect -50 207081 50 207097
rect -50 207023 50 207039
rect -50 206989 -34 207023
rect 34 206989 50 207023
rect -50 206951 50 206989
rect -50 205913 50 205951
rect -50 205879 -34 205913
rect 34 205879 50 205913
rect -50 205863 50 205879
rect -50 205805 50 205821
rect -50 205771 -34 205805
rect 34 205771 50 205805
rect -50 205733 50 205771
rect -50 204695 50 204733
rect -50 204661 -34 204695
rect 34 204661 50 204695
rect -50 204645 50 204661
rect -50 204587 50 204603
rect -50 204553 -34 204587
rect 34 204553 50 204587
rect -50 204515 50 204553
rect -50 203477 50 203515
rect -50 203443 -34 203477
rect 34 203443 50 203477
rect -50 203427 50 203443
rect -50 203369 50 203385
rect -50 203335 -34 203369
rect 34 203335 50 203369
rect -50 203297 50 203335
rect -50 202259 50 202297
rect -50 202225 -34 202259
rect 34 202225 50 202259
rect -50 202209 50 202225
rect -50 202151 50 202167
rect -50 202117 -34 202151
rect 34 202117 50 202151
rect -50 202079 50 202117
rect -50 201041 50 201079
rect -50 201007 -34 201041
rect 34 201007 50 201041
rect -50 200991 50 201007
rect -50 200933 50 200949
rect -50 200899 -34 200933
rect 34 200899 50 200933
rect -50 200861 50 200899
rect -50 199823 50 199861
rect -50 199789 -34 199823
rect 34 199789 50 199823
rect -50 199773 50 199789
rect -50 199715 50 199731
rect -50 199681 -34 199715
rect 34 199681 50 199715
rect -50 199643 50 199681
rect -50 198605 50 198643
rect -50 198571 -34 198605
rect 34 198571 50 198605
rect -50 198555 50 198571
rect -50 198497 50 198513
rect -50 198463 -34 198497
rect 34 198463 50 198497
rect -50 198425 50 198463
rect -50 197387 50 197425
rect -50 197353 -34 197387
rect 34 197353 50 197387
rect -50 197337 50 197353
rect -50 197279 50 197295
rect -50 197245 -34 197279
rect 34 197245 50 197279
rect -50 197207 50 197245
rect -50 196169 50 196207
rect -50 196135 -34 196169
rect 34 196135 50 196169
rect -50 196119 50 196135
rect -50 196061 50 196077
rect -50 196027 -34 196061
rect 34 196027 50 196061
rect -50 195989 50 196027
rect -50 194951 50 194989
rect -50 194917 -34 194951
rect 34 194917 50 194951
rect -50 194901 50 194917
rect -50 194843 50 194859
rect -50 194809 -34 194843
rect 34 194809 50 194843
rect -50 194771 50 194809
rect -50 193733 50 193771
rect -50 193699 -34 193733
rect 34 193699 50 193733
rect -50 193683 50 193699
rect -50 193625 50 193641
rect -50 193591 -34 193625
rect 34 193591 50 193625
rect -50 193553 50 193591
rect -50 192515 50 192553
rect -50 192481 -34 192515
rect 34 192481 50 192515
rect -50 192465 50 192481
rect -50 192407 50 192423
rect -50 192373 -34 192407
rect 34 192373 50 192407
rect -50 192335 50 192373
rect -50 191297 50 191335
rect -50 191263 -34 191297
rect 34 191263 50 191297
rect -50 191247 50 191263
rect -50 191189 50 191205
rect -50 191155 -34 191189
rect 34 191155 50 191189
rect -50 191117 50 191155
rect -50 190079 50 190117
rect -50 190045 -34 190079
rect 34 190045 50 190079
rect -50 190029 50 190045
rect -50 189971 50 189987
rect -50 189937 -34 189971
rect 34 189937 50 189971
rect -50 189899 50 189937
rect -50 188861 50 188899
rect -50 188827 -34 188861
rect 34 188827 50 188861
rect -50 188811 50 188827
rect -50 188753 50 188769
rect -50 188719 -34 188753
rect 34 188719 50 188753
rect -50 188681 50 188719
rect -50 187643 50 187681
rect -50 187609 -34 187643
rect 34 187609 50 187643
rect -50 187593 50 187609
rect -50 187535 50 187551
rect -50 187501 -34 187535
rect 34 187501 50 187535
rect -50 187463 50 187501
rect -50 186425 50 186463
rect -50 186391 -34 186425
rect 34 186391 50 186425
rect -50 186375 50 186391
rect -50 186317 50 186333
rect -50 186283 -34 186317
rect 34 186283 50 186317
rect -50 186245 50 186283
rect -50 185207 50 185245
rect -50 185173 -34 185207
rect 34 185173 50 185207
rect -50 185157 50 185173
rect -50 185099 50 185115
rect -50 185065 -34 185099
rect 34 185065 50 185099
rect -50 185027 50 185065
rect -50 183989 50 184027
rect -50 183955 -34 183989
rect 34 183955 50 183989
rect -50 183939 50 183955
rect -50 183881 50 183897
rect -50 183847 -34 183881
rect 34 183847 50 183881
rect -50 183809 50 183847
rect -50 182771 50 182809
rect -50 182737 -34 182771
rect 34 182737 50 182771
rect -50 182721 50 182737
rect -50 182663 50 182679
rect -50 182629 -34 182663
rect 34 182629 50 182663
rect -50 182591 50 182629
rect -50 181553 50 181591
rect -50 181519 -34 181553
rect 34 181519 50 181553
rect -50 181503 50 181519
rect -50 181445 50 181461
rect -50 181411 -34 181445
rect 34 181411 50 181445
rect -50 181373 50 181411
rect -50 180335 50 180373
rect -50 180301 -34 180335
rect 34 180301 50 180335
rect -50 180285 50 180301
rect -50 180227 50 180243
rect -50 180193 -34 180227
rect 34 180193 50 180227
rect -50 180155 50 180193
rect -50 179117 50 179155
rect -50 179083 -34 179117
rect 34 179083 50 179117
rect -50 179067 50 179083
rect -50 179009 50 179025
rect -50 178975 -34 179009
rect 34 178975 50 179009
rect -50 178937 50 178975
rect -50 177899 50 177937
rect -50 177865 -34 177899
rect 34 177865 50 177899
rect -50 177849 50 177865
rect -50 177791 50 177807
rect -50 177757 -34 177791
rect 34 177757 50 177791
rect -50 177719 50 177757
rect -50 176681 50 176719
rect -50 176647 -34 176681
rect 34 176647 50 176681
rect -50 176631 50 176647
rect -50 176573 50 176589
rect -50 176539 -34 176573
rect 34 176539 50 176573
rect -50 176501 50 176539
rect -50 175463 50 175501
rect -50 175429 -34 175463
rect 34 175429 50 175463
rect -50 175413 50 175429
rect -50 175355 50 175371
rect -50 175321 -34 175355
rect 34 175321 50 175355
rect -50 175283 50 175321
rect -50 174245 50 174283
rect -50 174211 -34 174245
rect 34 174211 50 174245
rect -50 174195 50 174211
rect -50 174137 50 174153
rect -50 174103 -34 174137
rect 34 174103 50 174137
rect -50 174065 50 174103
rect -50 173027 50 173065
rect -50 172993 -34 173027
rect 34 172993 50 173027
rect -50 172977 50 172993
rect -50 172919 50 172935
rect -50 172885 -34 172919
rect 34 172885 50 172919
rect -50 172847 50 172885
rect -50 171809 50 171847
rect -50 171775 -34 171809
rect 34 171775 50 171809
rect -50 171759 50 171775
rect -50 171701 50 171717
rect -50 171667 -34 171701
rect 34 171667 50 171701
rect -50 171629 50 171667
rect -50 170591 50 170629
rect -50 170557 -34 170591
rect 34 170557 50 170591
rect -50 170541 50 170557
rect -50 170483 50 170499
rect -50 170449 -34 170483
rect 34 170449 50 170483
rect -50 170411 50 170449
rect -50 169373 50 169411
rect -50 169339 -34 169373
rect 34 169339 50 169373
rect -50 169323 50 169339
rect -50 169265 50 169281
rect -50 169231 -34 169265
rect 34 169231 50 169265
rect -50 169193 50 169231
rect -50 168155 50 168193
rect -50 168121 -34 168155
rect 34 168121 50 168155
rect -50 168105 50 168121
rect -50 168047 50 168063
rect -50 168013 -34 168047
rect 34 168013 50 168047
rect -50 167975 50 168013
rect -50 166937 50 166975
rect -50 166903 -34 166937
rect 34 166903 50 166937
rect -50 166887 50 166903
rect -50 166829 50 166845
rect -50 166795 -34 166829
rect 34 166795 50 166829
rect -50 166757 50 166795
rect -50 165719 50 165757
rect -50 165685 -34 165719
rect 34 165685 50 165719
rect -50 165669 50 165685
rect -50 165611 50 165627
rect -50 165577 -34 165611
rect 34 165577 50 165611
rect -50 165539 50 165577
rect -50 164501 50 164539
rect -50 164467 -34 164501
rect 34 164467 50 164501
rect -50 164451 50 164467
rect -50 164393 50 164409
rect -50 164359 -34 164393
rect 34 164359 50 164393
rect -50 164321 50 164359
rect -50 163283 50 163321
rect -50 163249 -34 163283
rect 34 163249 50 163283
rect -50 163233 50 163249
rect -50 163175 50 163191
rect -50 163141 -34 163175
rect 34 163141 50 163175
rect -50 163103 50 163141
rect -50 162065 50 162103
rect -50 162031 -34 162065
rect 34 162031 50 162065
rect -50 162015 50 162031
rect -50 161957 50 161973
rect -50 161923 -34 161957
rect 34 161923 50 161957
rect -50 161885 50 161923
rect -50 160847 50 160885
rect -50 160813 -34 160847
rect 34 160813 50 160847
rect -50 160797 50 160813
rect -50 160739 50 160755
rect -50 160705 -34 160739
rect 34 160705 50 160739
rect -50 160667 50 160705
rect -50 159629 50 159667
rect -50 159595 -34 159629
rect 34 159595 50 159629
rect -50 159579 50 159595
rect -50 159521 50 159537
rect -50 159487 -34 159521
rect 34 159487 50 159521
rect -50 159449 50 159487
rect -50 158411 50 158449
rect -50 158377 -34 158411
rect 34 158377 50 158411
rect -50 158361 50 158377
rect -50 158303 50 158319
rect -50 158269 -34 158303
rect 34 158269 50 158303
rect -50 158231 50 158269
rect -50 157193 50 157231
rect -50 157159 -34 157193
rect 34 157159 50 157193
rect -50 157143 50 157159
rect -50 157085 50 157101
rect -50 157051 -34 157085
rect 34 157051 50 157085
rect -50 157013 50 157051
rect -50 155975 50 156013
rect -50 155941 -34 155975
rect 34 155941 50 155975
rect -50 155925 50 155941
rect -50 155867 50 155883
rect -50 155833 -34 155867
rect 34 155833 50 155867
rect -50 155795 50 155833
rect -50 154757 50 154795
rect -50 154723 -34 154757
rect 34 154723 50 154757
rect -50 154707 50 154723
rect -50 154649 50 154665
rect -50 154615 -34 154649
rect 34 154615 50 154649
rect -50 154577 50 154615
rect -50 153539 50 153577
rect -50 153505 -34 153539
rect 34 153505 50 153539
rect -50 153489 50 153505
rect -50 153431 50 153447
rect -50 153397 -34 153431
rect 34 153397 50 153431
rect -50 153359 50 153397
rect -50 152321 50 152359
rect -50 152287 -34 152321
rect 34 152287 50 152321
rect -50 152271 50 152287
rect -50 152213 50 152229
rect -50 152179 -34 152213
rect 34 152179 50 152213
rect -50 152141 50 152179
rect -50 151103 50 151141
rect -50 151069 -34 151103
rect 34 151069 50 151103
rect -50 151053 50 151069
rect -50 150995 50 151011
rect -50 150961 -34 150995
rect 34 150961 50 150995
rect -50 150923 50 150961
rect -50 149885 50 149923
rect -50 149851 -34 149885
rect 34 149851 50 149885
rect -50 149835 50 149851
rect -50 149777 50 149793
rect -50 149743 -34 149777
rect 34 149743 50 149777
rect -50 149705 50 149743
rect -50 148667 50 148705
rect -50 148633 -34 148667
rect 34 148633 50 148667
rect -50 148617 50 148633
rect -50 148559 50 148575
rect -50 148525 -34 148559
rect 34 148525 50 148559
rect -50 148487 50 148525
rect -50 147449 50 147487
rect -50 147415 -34 147449
rect 34 147415 50 147449
rect -50 147399 50 147415
rect -50 147341 50 147357
rect -50 147307 -34 147341
rect 34 147307 50 147341
rect -50 147269 50 147307
rect -50 146231 50 146269
rect -50 146197 -34 146231
rect 34 146197 50 146231
rect -50 146181 50 146197
rect -50 146123 50 146139
rect -50 146089 -34 146123
rect 34 146089 50 146123
rect -50 146051 50 146089
rect -50 145013 50 145051
rect -50 144979 -34 145013
rect 34 144979 50 145013
rect -50 144963 50 144979
rect -50 144905 50 144921
rect -50 144871 -34 144905
rect 34 144871 50 144905
rect -50 144833 50 144871
rect -50 143795 50 143833
rect -50 143761 -34 143795
rect 34 143761 50 143795
rect -50 143745 50 143761
rect -50 143687 50 143703
rect -50 143653 -34 143687
rect 34 143653 50 143687
rect -50 143615 50 143653
rect -50 142577 50 142615
rect -50 142543 -34 142577
rect 34 142543 50 142577
rect -50 142527 50 142543
rect -50 142469 50 142485
rect -50 142435 -34 142469
rect 34 142435 50 142469
rect -50 142397 50 142435
rect -50 141359 50 141397
rect -50 141325 -34 141359
rect 34 141325 50 141359
rect -50 141309 50 141325
rect -50 141251 50 141267
rect -50 141217 -34 141251
rect 34 141217 50 141251
rect -50 141179 50 141217
rect -50 140141 50 140179
rect -50 140107 -34 140141
rect 34 140107 50 140141
rect -50 140091 50 140107
rect -50 140033 50 140049
rect -50 139999 -34 140033
rect 34 139999 50 140033
rect -50 139961 50 139999
rect -50 138923 50 138961
rect -50 138889 -34 138923
rect 34 138889 50 138923
rect -50 138873 50 138889
rect -50 138815 50 138831
rect -50 138781 -34 138815
rect 34 138781 50 138815
rect -50 138743 50 138781
rect -50 137705 50 137743
rect -50 137671 -34 137705
rect 34 137671 50 137705
rect -50 137655 50 137671
rect -50 137597 50 137613
rect -50 137563 -34 137597
rect 34 137563 50 137597
rect -50 137525 50 137563
rect -50 136487 50 136525
rect -50 136453 -34 136487
rect 34 136453 50 136487
rect -50 136437 50 136453
rect -50 136379 50 136395
rect -50 136345 -34 136379
rect 34 136345 50 136379
rect -50 136307 50 136345
rect -50 135269 50 135307
rect -50 135235 -34 135269
rect 34 135235 50 135269
rect -50 135219 50 135235
rect -50 135161 50 135177
rect -50 135127 -34 135161
rect 34 135127 50 135161
rect -50 135089 50 135127
rect -50 134051 50 134089
rect -50 134017 -34 134051
rect 34 134017 50 134051
rect -50 134001 50 134017
rect -50 133943 50 133959
rect -50 133909 -34 133943
rect 34 133909 50 133943
rect -50 133871 50 133909
rect -50 132833 50 132871
rect -50 132799 -34 132833
rect 34 132799 50 132833
rect -50 132783 50 132799
rect -50 132725 50 132741
rect -50 132691 -34 132725
rect 34 132691 50 132725
rect -50 132653 50 132691
rect -50 131615 50 131653
rect -50 131581 -34 131615
rect 34 131581 50 131615
rect -50 131565 50 131581
rect -50 131507 50 131523
rect -50 131473 -34 131507
rect 34 131473 50 131507
rect -50 131435 50 131473
rect -50 130397 50 130435
rect -50 130363 -34 130397
rect 34 130363 50 130397
rect -50 130347 50 130363
rect -50 130289 50 130305
rect -50 130255 -34 130289
rect 34 130255 50 130289
rect -50 130217 50 130255
rect -50 129179 50 129217
rect -50 129145 -34 129179
rect 34 129145 50 129179
rect -50 129129 50 129145
rect -50 129071 50 129087
rect -50 129037 -34 129071
rect 34 129037 50 129071
rect -50 128999 50 129037
rect -50 127961 50 127999
rect -50 127927 -34 127961
rect 34 127927 50 127961
rect -50 127911 50 127927
rect -50 127853 50 127869
rect -50 127819 -34 127853
rect 34 127819 50 127853
rect -50 127781 50 127819
rect -50 126743 50 126781
rect -50 126709 -34 126743
rect 34 126709 50 126743
rect -50 126693 50 126709
rect -50 126635 50 126651
rect -50 126601 -34 126635
rect 34 126601 50 126635
rect -50 126563 50 126601
rect -50 125525 50 125563
rect -50 125491 -34 125525
rect 34 125491 50 125525
rect -50 125475 50 125491
rect -50 125417 50 125433
rect -50 125383 -34 125417
rect 34 125383 50 125417
rect -50 125345 50 125383
rect -50 124307 50 124345
rect -50 124273 -34 124307
rect 34 124273 50 124307
rect -50 124257 50 124273
rect -50 124199 50 124215
rect -50 124165 -34 124199
rect 34 124165 50 124199
rect -50 124127 50 124165
rect -50 123089 50 123127
rect -50 123055 -34 123089
rect 34 123055 50 123089
rect -50 123039 50 123055
rect -50 122981 50 122997
rect -50 122947 -34 122981
rect 34 122947 50 122981
rect -50 122909 50 122947
rect -50 121871 50 121909
rect -50 121837 -34 121871
rect 34 121837 50 121871
rect -50 121821 50 121837
rect -50 121763 50 121779
rect -50 121729 -34 121763
rect 34 121729 50 121763
rect -50 121691 50 121729
rect -50 120653 50 120691
rect -50 120619 -34 120653
rect 34 120619 50 120653
rect -50 120603 50 120619
rect -50 120545 50 120561
rect -50 120511 -34 120545
rect 34 120511 50 120545
rect -50 120473 50 120511
rect -50 119435 50 119473
rect -50 119401 -34 119435
rect 34 119401 50 119435
rect -50 119385 50 119401
rect -50 119327 50 119343
rect -50 119293 -34 119327
rect 34 119293 50 119327
rect -50 119255 50 119293
rect -50 118217 50 118255
rect -50 118183 -34 118217
rect 34 118183 50 118217
rect -50 118167 50 118183
rect -50 118109 50 118125
rect -50 118075 -34 118109
rect 34 118075 50 118109
rect -50 118037 50 118075
rect -50 116999 50 117037
rect -50 116965 -34 116999
rect 34 116965 50 116999
rect -50 116949 50 116965
rect -50 116891 50 116907
rect -50 116857 -34 116891
rect 34 116857 50 116891
rect -50 116819 50 116857
rect -50 115781 50 115819
rect -50 115747 -34 115781
rect 34 115747 50 115781
rect -50 115731 50 115747
rect -50 115673 50 115689
rect -50 115639 -34 115673
rect 34 115639 50 115673
rect -50 115601 50 115639
rect -50 114563 50 114601
rect -50 114529 -34 114563
rect 34 114529 50 114563
rect -50 114513 50 114529
rect -50 114455 50 114471
rect -50 114421 -34 114455
rect 34 114421 50 114455
rect -50 114383 50 114421
rect -50 113345 50 113383
rect -50 113311 -34 113345
rect 34 113311 50 113345
rect -50 113295 50 113311
rect -50 113237 50 113253
rect -50 113203 -34 113237
rect 34 113203 50 113237
rect -50 113165 50 113203
rect -50 112127 50 112165
rect -50 112093 -34 112127
rect 34 112093 50 112127
rect -50 112077 50 112093
rect -50 112019 50 112035
rect -50 111985 -34 112019
rect 34 111985 50 112019
rect -50 111947 50 111985
rect -50 110909 50 110947
rect -50 110875 -34 110909
rect 34 110875 50 110909
rect -50 110859 50 110875
rect -50 110801 50 110817
rect -50 110767 -34 110801
rect 34 110767 50 110801
rect -50 110729 50 110767
rect -50 109691 50 109729
rect -50 109657 -34 109691
rect 34 109657 50 109691
rect -50 109641 50 109657
rect -50 109583 50 109599
rect -50 109549 -34 109583
rect 34 109549 50 109583
rect -50 109511 50 109549
rect -50 108473 50 108511
rect -50 108439 -34 108473
rect 34 108439 50 108473
rect -50 108423 50 108439
rect -50 108365 50 108381
rect -50 108331 -34 108365
rect 34 108331 50 108365
rect -50 108293 50 108331
rect -50 107255 50 107293
rect -50 107221 -34 107255
rect 34 107221 50 107255
rect -50 107205 50 107221
rect -50 107147 50 107163
rect -50 107113 -34 107147
rect 34 107113 50 107147
rect -50 107075 50 107113
rect -50 106037 50 106075
rect -50 106003 -34 106037
rect 34 106003 50 106037
rect -50 105987 50 106003
rect -50 105929 50 105945
rect -50 105895 -34 105929
rect 34 105895 50 105929
rect -50 105857 50 105895
rect -50 104819 50 104857
rect -50 104785 -34 104819
rect 34 104785 50 104819
rect -50 104769 50 104785
rect -50 104711 50 104727
rect -50 104677 -34 104711
rect 34 104677 50 104711
rect -50 104639 50 104677
rect -50 103601 50 103639
rect -50 103567 -34 103601
rect 34 103567 50 103601
rect -50 103551 50 103567
rect -50 103493 50 103509
rect -50 103459 -34 103493
rect 34 103459 50 103493
rect -50 103421 50 103459
rect -50 102383 50 102421
rect -50 102349 -34 102383
rect 34 102349 50 102383
rect -50 102333 50 102349
rect -50 102275 50 102291
rect -50 102241 -34 102275
rect 34 102241 50 102275
rect -50 102203 50 102241
rect -50 101165 50 101203
rect -50 101131 -34 101165
rect 34 101131 50 101165
rect -50 101115 50 101131
rect -50 101057 50 101073
rect -50 101023 -34 101057
rect 34 101023 50 101057
rect -50 100985 50 101023
rect -50 99947 50 99985
rect -50 99913 -34 99947
rect 34 99913 50 99947
rect -50 99897 50 99913
rect -50 99839 50 99855
rect -50 99805 -34 99839
rect 34 99805 50 99839
rect -50 99767 50 99805
rect -50 98729 50 98767
rect -50 98695 -34 98729
rect 34 98695 50 98729
rect -50 98679 50 98695
rect -50 98621 50 98637
rect -50 98587 -34 98621
rect 34 98587 50 98621
rect -50 98549 50 98587
rect -50 97511 50 97549
rect -50 97477 -34 97511
rect 34 97477 50 97511
rect -50 97461 50 97477
rect -50 97403 50 97419
rect -50 97369 -34 97403
rect 34 97369 50 97403
rect -50 97331 50 97369
rect -50 96293 50 96331
rect -50 96259 -34 96293
rect 34 96259 50 96293
rect -50 96243 50 96259
rect -50 96185 50 96201
rect -50 96151 -34 96185
rect 34 96151 50 96185
rect -50 96113 50 96151
rect -50 95075 50 95113
rect -50 95041 -34 95075
rect 34 95041 50 95075
rect -50 95025 50 95041
rect -50 94967 50 94983
rect -50 94933 -34 94967
rect 34 94933 50 94967
rect -50 94895 50 94933
rect -50 93857 50 93895
rect -50 93823 -34 93857
rect 34 93823 50 93857
rect -50 93807 50 93823
rect -50 93749 50 93765
rect -50 93715 -34 93749
rect 34 93715 50 93749
rect -50 93677 50 93715
rect -50 92639 50 92677
rect -50 92605 -34 92639
rect 34 92605 50 92639
rect -50 92589 50 92605
rect -50 92531 50 92547
rect -50 92497 -34 92531
rect 34 92497 50 92531
rect -50 92459 50 92497
rect -50 91421 50 91459
rect -50 91387 -34 91421
rect 34 91387 50 91421
rect -50 91371 50 91387
rect -50 91313 50 91329
rect -50 91279 -34 91313
rect 34 91279 50 91313
rect -50 91241 50 91279
rect -50 90203 50 90241
rect -50 90169 -34 90203
rect 34 90169 50 90203
rect -50 90153 50 90169
rect -50 90095 50 90111
rect -50 90061 -34 90095
rect 34 90061 50 90095
rect -50 90023 50 90061
rect -50 88985 50 89023
rect -50 88951 -34 88985
rect 34 88951 50 88985
rect -50 88935 50 88951
rect -50 88877 50 88893
rect -50 88843 -34 88877
rect 34 88843 50 88877
rect -50 88805 50 88843
rect -50 87767 50 87805
rect -50 87733 -34 87767
rect 34 87733 50 87767
rect -50 87717 50 87733
rect -50 87659 50 87675
rect -50 87625 -34 87659
rect 34 87625 50 87659
rect -50 87587 50 87625
rect -50 86549 50 86587
rect -50 86515 -34 86549
rect 34 86515 50 86549
rect -50 86499 50 86515
rect -50 86441 50 86457
rect -50 86407 -34 86441
rect 34 86407 50 86441
rect -50 86369 50 86407
rect -50 85331 50 85369
rect -50 85297 -34 85331
rect 34 85297 50 85331
rect -50 85281 50 85297
rect -50 85223 50 85239
rect -50 85189 -34 85223
rect 34 85189 50 85223
rect -50 85151 50 85189
rect -50 84113 50 84151
rect -50 84079 -34 84113
rect 34 84079 50 84113
rect -50 84063 50 84079
rect -50 84005 50 84021
rect -50 83971 -34 84005
rect 34 83971 50 84005
rect -50 83933 50 83971
rect -50 82895 50 82933
rect -50 82861 -34 82895
rect 34 82861 50 82895
rect -50 82845 50 82861
rect -50 82787 50 82803
rect -50 82753 -34 82787
rect 34 82753 50 82787
rect -50 82715 50 82753
rect -50 81677 50 81715
rect -50 81643 -34 81677
rect 34 81643 50 81677
rect -50 81627 50 81643
rect -50 81569 50 81585
rect -50 81535 -34 81569
rect 34 81535 50 81569
rect -50 81497 50 81535
rect -50 80459 50 80497
rect -50 80425 -34 80459
rect 34 80425 50 80459
rect -50 80409 50 80425
rect -50 80351 50 80367
rect -50 80317 -34 80351
rect 34 80317 50 80351
rect -50 80279 50 80317
rect -50 79241 50 79279
rect -50 79207 -34 79241
rect 34 79207 50 79241
rect -50 79191 50 79207
rect -50 79133 50 79149
rect -50 79099 -34 79133
rect 34 79099 50 79133
rect -50 79061 50 79099
rect -50 78023 50 78061
rect -50 77989 -34 78023
rect 34 77989 50 78023
rect -50 77973 50 77989
rect -50 77915 50 77931
rect -50 77881 -34 77915
rect 34 77881 50 77915
rect -50 77843 50 77881
rect -50 76805 50 76843
rect -50 76771 -34 76805
rect 34 76771 50 76805
rect -50 76755 50 76771
rect -50 76697 50 76713
rect -50 76663 -34 76697
rect 34 76663 50 76697
rect -50 76625 50 76663
rect -50 75587 50 75625
rect -50 75553 -34 75587
rect 34 75553 50 75587
rect -50 75537 50 75553
rect -50 75479 50 75495
rect -50 75445 -34 75479
rect 34 75445 50 75479
rect -50 75407 50 75445
rect -50 74369 50 74407
rect -50 74335 -34 74369
rect 34 74335 50 74369
rect -50 74319 50 74335
rect -50 74261 50 74277
rect -50 74227 -34 74261
rect 34 74227 50 74261
rect -50 74189 50 74227
rect -50 73151 50 73189
rect -50 73117 -34 73151
rect 34 73117 50 73151
rect -50 73101 50 73117
rect -50 73043 50 73059
rect -50 73009 -34 73043
rect 34 73009 50 73043
rect -50 72971 50 73009
rect -50 71933 50 71971
rect -50 71899 -34 71933
rect 34 71899 50 71933
rect -50 71883 50 71899
rect -50 71825 50 71841
rect -50 71791 -34 71825
rect 34 71791 50 71825
rect -50 71753 50 71791
rect -50 70715 50 70753
rect -50 70681 -34 70715
rect 34 70681 50 70715
rect -50 70665 50 70681
rect -50 70607 50 70623
rect -50 70573 -34 70607
rect 34 70573 50 70607
rect -50 70535 50 70573
rect -50 69497 50 69535
rect -50 69463 -34 69497
rect 34 69463 50 69497
rect -50 69447 50 69463
rect -50 69389 50 69405
rect -50 69355 -34 69389
rect 34 69355 50 69389
rect -50 69317 50 69355
rect -50 68279 50 68317
rect -50 68245 -34 68279
rect 34 68245 50 68279
rect -50 68229 50 68245
rect -50 68171 50 68187
rect -50 68137 -34 68171
rect 34 68137 50 68171
rect -50 68099 50 68137
rect -50 67061 50 67099
rect -50 67027 -34 67061
rect 34 67027 50 67061
rect -50 67011 50 67027
rect -50 66953 50 66969
rect -50 66919 -34 66953
rect 34 66919 50 66953
rect -50 66881 50 66919
rect -50 65843 50 65881
rect -50 65809 -34 65843
rect 34 65809 50 65843
rect -50 65793 50 65809
rect -50 65735 50 65751
rect -50 65701 -34 65735
rect 34 65701 50 65735
rect -50 65663 50 65701
rect -50 64625 50 64663
rect -50 64591 -34 64625
rect 34 64591 50 64625
rect -50 64575 50 64591
rect -50 64517 50 64533
rect -50 64483 -34 64517
rect 34 64483 50 64517
rect -50 64445 50 64483
rect -50 63407 50 63445
rect -50 63373 -34 63407
rect 34 63373 50 63407
rect -50 63357 50 63373
rect -50 63299 50 63315
rect -50 63265 -34 63299
rect 34 63265 50 63299
rect -50 63227 50 63265
rect -50 62189 50 62227
rect -50 62155 -34 62189
rect 34 62155 50 62189
rect -50 62139 50 62155
rect -50 62081 50 62097
rect -50 62047 -34 62081
rect 34 62047 50 62081
rect -50 62009 50 62047
rect -50 60971 50 61009
rect -50 60937 -34 60971
rect 34 60937 50 60971
rect -50 60921 50 60937
rect -50 60863 50 60879
rect -50 60829 -34 60863
rect 34 60829 50 60863
rect -50 60791 50 60829
rect -50 59753 50 59791
rect -50 59719 -34 59753
rect 34 59719 50 59753
rect -50 59703 50 59719
rect -50 59645 50 59661
rect -50 59611 -34 59645
rect 34 59611 50 59645
rect -50 59573 50 59611
rect -50 58535 50 58573
rect -50 58501 -34 58535
rect 34 58501 50 58535
rect -50 58485 50 58501
rect -50 58427 50 58443
rect -50 58393 -34 58427
rect 34 58393 50 58427
rect -50 58355 50 58393
rect -50 57317 50 57355
rect -50 57283 -34 57317
rect 34 57283 50 57317
rect -50 57267 50 57283
rect -50 57209 50 57225
rect -50 57175 -34 57209
rect 34 57175 50 57209
rect -50 57137 50 57175
rect -50 56099 50 56137
rect -50 56065 -34 56099
rect 34 56065 50 56099
rect -50 56049 50 56065
rect -50 55991 50 56007
rect -50 55957 -34 55991
rect 34 55957 50 55991
rect -50 55919 50 55957
rect -50 54881 50 54919
rect -50 54847 -34 54881
rect 34 54847 50 54881
rect -50 54831 50 54847
rect -50 54773 50 54789
rect -50 54739 -34 54773
rect 34 54739 50 54773
rect -50 54701 50 54739
rect -50 53663 50 53701
rect -50 53629 -34 53663
rect 34 53629 50 53663
rect -50 53613 50 53629
rect -50 53555 50 53571
rect -50 53521 -34 53555
rect 34 53521 50 53555
rect -50 53483 50 53521
rect -50 52445 50 52483
rect -50 52411 -34 52445
rect 34 52411 50 52445
rect -50 52395 50 52411
rect -50 52337 50 52353
rect -50 52303 -34 52337
rect 34 52303 50 52337
rect -50 52265 50 52303
rect -50 51227 50 51265
rect -50 51193 -34 51227
rect 34 51193 50 51227
rect -50 51177 50 51193
rect -50 51119 50 51135
rect -50 51085 -34 51119
rect 34 51085 50 51119
rect -50 51047 50 51085
rect -50 50009 50 50047
rect -50 49975 -34 50009
rect 34 49975 50 50009
rect -50 49959 50 49975
rect -50 49901 50 49917
rect -50 49867 -34 49901
rect 34 49867 50 49901
rect -50 49829 50 49867
rect -50 48791 50 48829
rect -50 48757 -34 48791
rect 34 48757 50 48791
rect -50 48741 50 48757
rect -50 48683 50 48699
rect -50 48649 -34 48683
rect 34 48649 50 48683
rect -50 48611 50 48649
rect -50 47573 50 47611
rect -50 47539 -34 47573
rect 34 47539 50 47573
rect -50 47523 50 47539
rect -50 47465 50 47481
rect -50 47431 -34 47465
rect 34 47431 50 47465
rect -50 47393 50 47431
rect -50 46355 50 46393
rect -50 46321 -34 46355
rect 34 46321 50 46355
rect -50 46305 50 46321
rect -50 46247 50 46263
rect -50 46213 -34 46247
rect 34 46213 50 46247
rect -50 46175 50 46213
rect -50 45137 50 45175
rect -50 45103 -34 45137
rect 34 45103 50 45137
rect -50 45087 50 45103
rect -50 45029 50 45045
rect -50 44995 -34 45029
rect 34 44995 50 45029
rect -50 44957 50 44995
rect -50 43919 50 43957
rect -50 43885 -34 43919
rect 34 43885 50 43919
rect -50 43869 50 43885
rect -50 43811 50 43827
rect -50 43777 -34 43811
rect 34 43777 50 43811
rect -50 43739 50 43777
rect -50 42701 50 42739
rect -50 42667 -34 42701
rect 34 42667 50 42701
rect -50 42651 50 42667
rect -50 42593 50 42609
rect -50 42559 -34 42593
rect 34 42559 50 42593
rect -50 42521 50 42559
rect -50 41483 50 41521
rect -50 41449 -34 41483
rect 34 41449 50 41483
rect -50 41433 50 41449
rect -50 41375 50 41391
rect -50 41341 -34 41375
rect 34 41341 50 41375
rect -50 41303 50 41341
rect -50 40265 50 40303
rect -50 40231 -34 40265
rect 34 40231 50 40265
rect -50 40215 50 40231
rect -50 40157 50 40173
rect -50 40123 -34 40157
rect 34 40123 50 40157
rect -50 40085 50 40123
rect -50 39047 50 39085
rect -50 39013 -34 39047
rect 34 39013 50 39047
rect -50 38997 50 39013
rect -50 38939 50 38955
rect -50 38905 -34 38939
rect 34 38905 50 38939
rect -50 38867 50 38905
rect -50 37829 50 37867
rect -50 37795 -34 37829
rect 34 37795 50 37829
rect -50 37779 50 37795
rect -50 37721 50 37737
rect -50 37687 -34 37721
rect 34 37687 50 37721
rect -50 37649 50 37687
rect -50 36611 50 36649
rect -50 36577 -34 36611
rect 34 36577 50 36611
rect -50 36561 50 36577
rect -50 36503 50 36519
rect -50 36469 -34 36503
rect 34 36469 50 36503
rect -50 36431 50 36469
rect -50 35393 50 35431
rect -50 35359 -34 35393
rect 34 35359 50 35393
rect -50 35343 50 35359
rect -50 35285 50 35301
rect -50 35251 -34 35285
rect 34 35251 50 35285
rect -50 35213 50 35251
rect -50 34175 50 34213
rect -50 34141 -34 34175
rect 34 34141 50 34175
rect -50 34125 50 34141
rect -50 34067 50 34083
rect -50 34033 -34 34067
rect 34 34033 50 34067
rect -50 33995 50 34033
rect -50 32957 50 32995
rect -50 32923 -34 32957
rect 34 32923 50 32957
rect -50 32907 50 32923
rect -50 32849 50 32865
rect -50 32815 -34 32849
rect 34 32815 50 32849
rect -50 32777 50 32815
rect -50 31739 50 31777
rect -50 31705 -34 31739
rect 34 31705 50 31739
rect -50 31689 50 31705
rect -50 31631 50 31647
rect -50 31597 -34 31631
rect 34 31597 50 31631
rect -50 31559 50 31597
rect -50 30521 50 30559
rect -50 30487 -34 30521
rect 34 30487 50 30521
rect -50 30471 50 30487
rect -50 30413 50 30429
rect -50 30379 -34 30413
rect 34 30379 50 30413
rect -50 30341 50 30379
rect -50 29303 50 29341
rect -50 29269 -34 29303
rect 34 29269 50 29303
rect -50 29253 50 29269
rect -50 29195 50 29211
rect -50 29161 -34 29195
rect 34 29161 50 29195
rect -50 29123 50 29161
rect -50 28085 50 28123
rect -50 28051 -34 28085
rect 34 28051 50 28085
rect -50 28035 50 28051
rect -50 27977 50 27993
rect -50 27943 -34 27977
rect 34 27943 50 27977
rect -50 27905 50 27943
rect -50 26867 50 26905
rect -50 26833 -34 26867
rect 34 26833 50 26867
rect -50 26817 50 26833
rect -50 26759 50 26775
rect -50 26725 -34 26759
rect 34 26725 50 26759
rect -50 26687 50 26725
rect -50 25649 50 25687
rect -50 25615 -34 25649
rect 34 25615 50 25649
rect -50 25599 50 25615
rect -50 25541 50 25557
rect -50 25507 -34 25541
rect 34 25507 50 25541
rect -50 25469 50 25507
rect -50 24431 50 24469
rect -50 24397 -34 24431
rect 34 24397 50 24431
rect -50 24381 50 24397
rect -50 24323 50 24339
rect -50 24289 -34 24323
rect 34 24289 50 24323
rect -50 24251 50 24289
rect -50 23213 50 23251
rect -50 23179 -34 23213
rect 34 23179 50 23213
rect -50 23163 50 23179
rect -50 23105 50 23121
rect -50 23071 -34 23105
rect 34 23071 50 23105
rect -50 23033 50 23071
rect -50 21995 50 22033
rect -50 21961 -34 21995
rect 34 21961 50 21995
rect -50 21945 50 21961
rect -50 21887 50 21903
rect -50 21853 -34 21887
rect 34 21853 50 21887
rect -50 21815 50 21853
rect -50 20777 50 20815
rect -50 20743 -34 20777
rect 34 20743 50 20777
rect -50 20727 50 20743
rect -50 20669 50 20685
rect -50 20635 -34 20669
rect 34 20635 50 20669
rect -50 20597 50 20635
rect -50 19559 50 19597
rect -50 19525 -34 19559
rect 34 19525 50 19559
rect -50 19509 50 19525
rect -50 19451 50 19467
rect -50 19417 -34 19451
rect 34 19417 50 19451
rect -50 19379 50 19417
rect -50 18341 50 18379
rect -50 18307 -34 18341
rect 34 18307 50 18341
rect -50 18291 50 18307
rect -50 18233 50 18249
rect -50 18199 -34 18233
rect 34 18199 50 18233
rect -50 18161 50 18199
rect -50 17123 50 17161
rect -50 17089 -34 17123
rect 34 17089 50 17123
rect -50 17073 50 17089
rect -50 17015 50 17031
rect -50 16981 -34 17015
rect 34 16981 50 17015
rect -50 16943 50 16981
rect -50 15905 50 15943
rect -50 15871 -34 15905
rect 34 15871 50 15905
rect -50 15855 50 15871
rect -50 15797 50 15813
rect -50 15763 -34 15797
rect 34 15763 50 15797
rect -50 15725 50 15763
rect -50 14687 50 14725
rect -50 14653 -34 14687
rect 34 14653 50 14687
rect -50 14637 50 14653
rect -50 14579 50 14595
rect -50 14545 -34 14579
rect 34 14545 50 14579
rect -50 14507 50 14545
rect -50 13469 50 13507
rect -50 13435 -34 13469
rect 34 13435 50 13469
rect -50 13419 50 13435
rect -50 13361 50 13377
rect -50 13327 -34 13361
rect 34 13327 50 13361
rect -50 13289 50 13327
rect -50 12251 50 12289
rect -50 12217 -34 12251
rect 34 12217 50 12251
rect -50 12201 50 12217
rect -50 12143 50 12159
rect -50 12109 -34 12143
rect 34 12109 50 12143
rect -50 12071 50 12109
rect -50 11033 50 11071
rect -50 10999 -34 11033
rect 34 10999 50 11033
rect -50 10983 50 10999
rect -50 10925 50 10941
rect -50 10891 -34 10925
rect 34 10891 50 10925
rect -50 10853 50 10891
rect -50 9815 50 9853
rect -50 9781 -34 9815
rect 34 9781 50 9815
rect -50 9765 50 9781
rect -50 9707 50 9723
rect -50 9673 -34 9707
rect 34 9673 50 9707
rect -50 9635 50 9673
rect -50 8597 50 8635
rect -50 8563 -34 8597
rect 34 8563 50 8597
rect -50 8547 50 8563
rect -50 8489 50 8505
rect -50 8455 -34 8489
rect 34 8455 50 8489
rect -50 8417 50 8455
rect -50 7379 50 7417
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -50 7329 50 7345
rect -50 7271 50 7287
rect -50 7237 -34 7271
rect 34 7237 50 7271
rect -50 7199 50 7237
rect -50 6161 50 6199
rect -50 6127 -34 6161
rect 34 6127 50 6161
rect -50 6111 50 6127
rect -50 6053 50 6069
rect -50 6019 -34 6053
rect 34 6019 50 6053
rect -50 5981 50 6019
rect -50 4943 50 4981
rect -50 4909 -34 4943
rect 34 4909 50 4943
rect -50 4893 50 4909
rect -50 4835 50 4851
rect -50 4801 -34 4835
rect 34 4801 50 4835
rect -50 4763 50 4801
rect -50 3725 50 3763
rect -50 3691 -34 3725
rect 34 3691 50 3725
rect -50 3675 50 3691
rect -50 3617 50 3633
rect -50 3583 -34 3617
rect 34 3583 50 3617
rect -50 3545 50 3583
rect -50 2507 50 2545
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -50 2457 50 2473
rect -50 2399 50 2415
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -50 2327 50 2365
rect -50 1289 50 1327
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1239 50 1255
rect -50 1181 50 1197
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -50 1109 50 1147
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -1147 50 -1109
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1197 50 -1181
rect -50 -1255 50 -1239
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -50 -1327 50 -1289
rect -50 -2365 50 -2327
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -50 -2415 50 -2399
rect -50 -2473 50 -2457
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -50 -2545 50 -2507
rect -50 -3583 50 -3545
rect -50 -3617 -34 -3583
rect 34 -3617 50 -3583
rect -50 -3633 50 -3617
rect -50 -3691 50 -3675
rect -50 -3725 -34 -3691
rect 34 -3725 50 -3691
rect -50 -3763 50 -3725
rect -50 -4801 50 -4763
rect -50 -4835 -34 -4801
rect 34 -4835 50 -4801
rect -50 -4851 50 -4835
rect -50 -4909 50 -4893
rect -50 -4943 -34 -4909
rect 34 -4943 50 -4909
rect -50 -4981 50 -4943
rect -50 -6019 50 -5981
rect -50 -6053 -34 -6019
rect 34 -6053 50 -6019
rect -50 -6069 50 -6053
rect -50 -6127 50 -6111
rect -50 -6161 -34 -6127
rect 34 -6161 50 -6127
rect -50 -6199 50 -6161
rect -50 -7237 50 -7199
rect -50 -7271 -34 -7237
rect 34 -7271 50 -7237
rect -50 -7287 50 -7271
rect -50 -7345 50 -7329
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -50 -7417 50 -7379
rect -50 -8455 50 -8417
rect -50 -8489 -34 -8455
rect 34 -8489 50 -8455
rect -50 -8505 50 -8489
rect -50 -8563 50 -8547
rect -50 -8597 -34 -8563
rect 34 -8597 50 -8563
rect -50 -8635 50 -8597
rect -50 -9673 50 -9635
rect -50 -9707 -34 -9673
rect 34 -9707 50 -9673
rect -50 -9723 50 -9707
rect -50 -9781 50 -9765
rect -50 -9815 -34 -9781
rect 34 -9815 50 -9781
rect -50 -9853 50 -9815
rect -50 -10891 50 -10853
rect -50 -10925 -34 -10891
rect 34 -10925 50 -10891
rect -50 -10941 50 -10925
rect -50 -10999 50 -10983
rect -50 -11033 -34 -10999
rect 34 -11033 50 -10999
rect -50 -11071 50 -11033
rect -50 -12109 50 -12071
rect -50 -12143 -34 -12109
rect 34 -12143 50 -12109
rect -50 -12159 50 -12143
rect -50 -12217 50 -12201
rect -50 -12251 -34 -12217
rect 34 -12251 50 -12217
rect -50 -12289 50 -12251
rect -50 -13327 50 -13289
rect -50 -13361 -34 -13327
rect 34 -13361 50 -13327
rect -50 -13377 50 -13361
rect -50 -13435 50 -13419
rect -50 -13469 -34 -13435
rect 34 -13469 50 -13435
rect -50 -13507 50 -13469
rect -50 -14545 50 -14507
rect -50 -14579 -34 -14545
rect 34 -14579 50 -14545
rect -50 -14595 50 -14579
rect -50 -14653 50 -14637
rect -50 -14687 -34 -14653
rect 34 -14687 50 -14653
rect -50 -14725 50 -14687
rect -50 -15763 50 -15725
rect -50 -15797 -34 -15763
rect 34 -15797 50 -15763
rect -50 -15813 50 -15797
rect -50 -15871 50 -15855
rect -50 -15905 -34 -15871
rect 34 -15905 50 -15871
rect -50 -15943 50 -15905
rect -50 -16981 50 -16943
rect -50 -17015 -34 -16981
rect 34 -17015 50 -16981
rect -50 -17031 50 -17015
rect -50 -17089 50 -17073
rect -50 -17123 -34 -17089
rect 34 -17123 50 -17089
rect -50 -17161 50 -17123
rect -50 -18199 50 -18161
rect -50 -18233 -34 -18199
rect 34 -18233 50 -18199
rect -50 -18249 50 -18233
rect -50 -18307 50 -18291
rect -50 -18341 -34 -18307
rect 34 -18341 50 -18307
rect -50 -18379 50 -18341
rect -50 -19417 50 -19379
rect -50 -19451 -34 -19417
rect 34 -19451 50 -19417
rect -50 -19467 50 -19451
rect -50 -19525 50 -19509
rect -50 -19559 -34 -19525
rect 34 -19559 50 -19525
rect -50 -19597 50 -19559
rect -50 -20635 50 -20597
rect -50 -20669 -34 -20635
rect 34 -20669 50 -20635
rect -50 -20685 50 -20669
rect -50 -20743 50 -20727
rect -50 -20777 -34 -20743
rect 34 -20777 50 -20743
rect -50 -20815 50 -20777
rect -50 -21853 50 -21815
rect -50 -21887 -34 -21853
rect 34 -21887 50 -21853
rect -50 -21903 50 -21887
rect -50 -21961 50 -21945
rect -50 -21995 -34 -21961
rect 34 -21995 50 -21961
rect -50 -22033 50 -21995
rect -50 -23071 50 -23033
rect -50 -23105 -34 -23071
rect 34 -23105 50 -23071
rect -50 -23121 50 -23105
rect -50 -23179 50 -23163
rect -50 -23213 -34 -23179
rect 34 -23213 50 -23179
rect -50 -23251 50 -23213
rect -50 -24289 50 -24251
rect -50 -24323 -34 -24289
rect 34 -24323 50 -24289
rect -50 -24339 50 -24323
rect -50 -24397 50 -24381
rect -50 -24431 -34 -24397
rect 34 -24431 50 -24397
rect -50 -24469 50 -24431
rect -50 -25507 50 -25469
rect -50 -25541 -34 -25507
rect 34 -25541 50 -25507
rect -50 -25557 50 -25541
rect -50 -25615 50 -25599
rect -50 -25649 -34 -25615
rect 34 -25649 50 -25615
rect -50 -25687 50 -25649
rect -50 -26725 50 -26687
rect -50 -26759 -34 -26725
rect 34 -26759 50 -26725
rect -50 -26775 50 -26759
rect -50 -26833 50 -26817
rect -50 -26867 -34 -26833
rect 34 -26867 50 -26833
rect -50 -26905 50 -26867
rect -50 -27943 50 -27905
rect -50 -27977 -34 -27943
rect 34 -27977 50 -27943
rect -50 -27993 50 -27977
rect -50 -28051 50 -28035
rect -50 -28085 -34 -28051
rect 34 -28085 50 -28051
rect -50 -28123 50 -28085
rect -50 -29161 50 -29123
rect -50 -29195 -34 -29161
rect 34 -29195 50 -29161
rect -50 -29211 50 -29195
rect -50 -29269 50 -29253
rect -50 -29303 -34 -29269
rect 34 -29303 50 -29269
rect -50 -29341 50 -29303
rect -50 -30379 50 -30341
rect -50 -30413 -34 -30379
rect 34 -30413 50 -30379
rect -50 -30429 50 -30413
rect -50 -30487 50 -30471
rect -50 -30521 -34 -30487
rect 34 -30521 50 -30487
rect -50 -30559 50 -30521
rect -50 -31597 50 -31559
rect -50 -31631 -34 -31597
rect 34 -31631 50 -31597
rect -50 -31647 50 -31631
rect -50 -31705 50 -31689
rect -50 -31739 -34 -31705
rect 34 -31739 50 -31705
rect -50 -31777 50 -31739
rect -50 -32815 50 -32777
rect -50 -32849 -34 -32815
rect 34 -32849 50 -32815
rect -50 -32865 50 -32849
rect -50 -32923 50 -32907
rect -50 -32957 -34 -32923
rect 34 -32957 50 -32923
rect -50 -32995 50 -32957
rect -50 -34033 50 -33995
rect -50 -34067 -34 -34033
rect 34 -34067 50 -34033
rect -50 -34083 50 -34067
rect -50 -34141 50 -34125
rect -50 -34175 -34 -34141
rect 34 -34175 50 -34141
rect -50 -34213 50 -34175
rect -50 -35251 50 -35213
rect -50 -35285 -34 -35251
rect 34 -35285 50 -35251
rect -50 -35301 50 -35285
rect -50 -35359 50 -35343
rect -50 -35393 -34 -35359
rect 34 -35393 50 -35359
rect -50 -35431 50 -35393
rect -50 -36469 50 -36431
rect -50 -36503 -34 -36469
rect 34 -36503 50 -36469
rect -50 -36519 50 -36503
rect -50 -36577 50 -36561
rect -50 -36611 -34 -36577
rect 34 -36611 50 -36577
rect -50 -36649 50 -36611
rect -50 -37687 50 -37649
rect -50 -37721 -34 -37687
rect 34 -37721 50 -37687
rect -50 -37737 50 -37721
rect -50 -37795 50 -37779
rect -50 -37829 -34 -37795
rect 34 -37829 50 -37795
rect -50 -37867 50 -37829
rect -50 -38905 50 -38867
rect -50 -38939 -34 -38905
rect 34 -38939 50 -38905
rect -50 -38955 50 -38939
rect -50 -39013 50 -38997
rect -50 -39047 -34 -39013
rect 34 -39047 50 -39013
rect -50 -39085 50 -39047
rect -50 -40123 50 -40085
rect -50 -40157 -34 -40123
rect 34 -40157 50 -40123
rect -50 -40173 50 -40157
rect -50 -40231 50 -40215
rect -50 -40265 -34 -40231
rect 34 -40265 50 -40231
rect -50 -40303 50 -40265
rect -50 -41341 50 -41303
rect -50 -41375 -34 -41341
rect 34 -41375 50 -41341
rect -50 -41391 50 -41375
rect -50 -41449 50 -41433
rect -50 -41483 -34 -41449
rect 34 -41483 50 -41449
rect -50 -41521 50 -41483
rect -50 -42559 50 -42521
rect -50 -42593 -34 -42559
rect 34 -42593 50 -42559
rect -50 -42609 50 -42593
rect -50 -42667 50 -42651
rect -50 -42701 -34 -42667
rect 34 -42701 50 -42667
rect -50 -42739 50 -42701
rect -50 -43777 50 -43739
rect -50 -43811 -34 -43777
rect 34 -43811 50 -43777
rect -50 -43827 50 -43811
rect -50 -43885 50 -43869
rect -50 -43919 -34 -43885
rect 34 -43919 50 -43885
rect -50 -43957 50 -43919
rect -50 -44995 50 -44957
rect -50 -45029 -34 -44995
rect 34 -45029 50 -44995
rect -50 -45045 50 -45029
rect -50 -45103 50 -45087
rect -50 -45137 -34 -45103
rect 34 -45137 50 -45103
rect -50 -45175 50 -45137
rect -50 -46213 50 -46175
rect -50 -46247 -34 -46213
rect 34 -46247 50 -46213
rect -50 -46263 50 -46247
rect -50 -46321 50 -46305
rect -50 -46355 -34 -46321
rect 34 -46355 50 -46321
rect -50 -46393 50 -46355
rect -50 -47431 50 -47393
rect -50 -47465 -34 -47431
rect 34 -47465 50 -47431
rect -50 -47481 50 -47465
rect -50 -47539 50 -47523
rect -50 -47573 -34 -47539
rect 34 -47573 50 -47539
rect -50 -47611 50 -47573
rect -50 -48649 50 -48611
rect -50 -48683 -34 -48649
rect 34 -48683 50 -48649
rect -50 -48699 50 -48683
rect -50 -48757 50 -48741
rect -50 -48791 -34 -48757
rect 34 -48791 50 -48757
rect -50 -48829 50 -48791
rect -50 -49867 50 -49829
rect -50 -49901 -34 -49867
rect 34 -49901 50 -49867
rect -50 -49917 50 -49901
rect -50 -49975 50 -49959
rect -50 -50009 -34 -49975
rect 34 -50009 50 -49975
rect -50 -50047 50 -50009
rect -50 -51085 50 -51047
rect -50 -51119 -34 -51085
rect 34 -51119 50 -51085
rect -50 -51135 50 -51119
rect -50 -51193 50 -51177
rect -50 -51227 -34 -51193
rect 34 -51227 50 -51193
rect -50 -51265 50 -51227
rect -50 -52303 50 -52265
rect -50 -52337 -34 -52303
rect 34 -52337 50 -52303
rect -50 -52353 50 -52337
rect -50 -52411 50 -52395
rect -50 -52445 -34 -52411
rect 34 -52445 50 -52411
rect -50 -52483 50 -52445
rect -50 -53521 50 -53483
rect -50 -53555 -34 -53521
rect 34 -53555 50 -53521
rect -50 -53571 50 -53555
rect -50 -53629 50 -53613
rect -50 -53663 -34 -53629
rect 34 -53663 50 -53629
rect -50 -53701 50 -53663
rect -50 -54739 50 -54701
rect -50 -54773 -34 -54739
rect 34 -54773 50 -54739
rect -50 -54789 50 -54773
rect -50 -54847 50 -54831
rect -50 -54881 -34 -54847
rect 34 -54881 50 -54847
rect -50 -54919 50 -54881
rect -50 -55957 50 -55919
rect -50 -55991 -34 -55957
rect 34 -55991 50 -55957
rect -50 -56007 50 -55991
rect -50 -56065 50 -56049
rect -50 -56099 -34 -56065
rect 34 -56099 50 -56065
rect -50 -56137 50 -56099
rect -50 -57175 50 -57137
rect -50 -57209 -34 -57175
rect 34 -57209 50 -57175
rect -50 -57225 50 -57209
rect -50 -57283 50 -57267
rect -50 -57317 -34 -57283
rect 34 -57317 50 -57283
rect -50 -57355 50 -57317
rect -50 -58393 50 -58355
rect -50 -58427 -34 -58393
rect 34 -58427 50 -58393
rect -50 -58443 50 -58427
rect -50 -58501 50 -58485
rect -50 -58535 -34 -58501
rect 34 -58535 50 -58501
rect -50 -58573 50 -58535
rect -50 -59611 50 -59573
rect -50 -59645 -34 -59611
rect 34 -59645 50 -59611
rect -50 -59661 50 -59645
rect -50 -59719 50 -59703
rect -50 -59753 -34 -59719
rect 34 -59753 50 -59719
rect -50 -59791 50 -59753
rect -50 -60829 50 -60791
rect -50 -60863 -34 -60829
rect 34 -60863 50 -60829
rect -50 -60879 50 -60863
rect -50 -60937 50 -60921
rect -50 -60971 -34 -60937
rect 34 -60971 50 -60937
rect -50 -61009 50 -60971
rect -50 -62047 50 -62009
rect -50 -62081 -34 -62047
rect 34 -62081 50 -62047
rect -50 -62097 50 -62081
rect -50 -62155 50 -62139
rect -50 -62189 -34 -62155
rect 34 -62189 50 -62155
rect -50 -62227 50 -62189
rect -50 -63265 50 -63227
rect -50 -63299 -34 -63265
rect 34 -63299 50 -63265
rect -50 -63315 50 -63299
rect -50 -63373 50 -63357
rect -50 -63407 -34 -63373
rect 34 -63407 50 -63373
rect -50 -63445 50 -63407
rect -50 -64483 50 -64445
rect -50 -64517 -34 -64483
rect 34 -64517 50 -64483
rect -50 -64533 50 -64517
rect -50 -64591 50 -64575
rect -50 -64625 -34 -64591
rect 34 -64625 50 -64591
rect -50 -64663 50 -64625
rect -50 -65701 50 -65663
rect -50 -65735 -34 -65701
rect 34 -65735 50 -65701
rect -50 -65751 50 -65735
rect -50 -65809 50 -65793
rect -50 -65843 -34 -65809
rect 34 -65843 50 -65809
rect -50 -65881 50 -65843
rect -50 -66919 50 -66881
rect -50 -66953 -34 -66919
rect 34 -66953 50 -66919
rect -50 -66969 50 -66953
rect -50 -67027 50 -67011
rect -50 -67061 -34 -67027
rect 34 -67061 50 -67027
rect -50 -67099 50 -67061
rect -50 -68137 50 -68099
rect -50 -68171 -34 -68137
rect 34 -68171 50 -68137
rect -50 -68187 50 -68171
rect -50 -68245 50 -68229
rect -50 -68279 -34 -68245
rect 34 -68279 50 -68245
rect -50 -68317 50 -68279
rect -50 -69355 50 -69317
rect -50 -69389 -34 -69355
rect 34 -69389 50 -69355
rect -50 -69405 50 -69389
rect -50 -69463 50 -69447
rect -50 -69497 -34 -69463
rect 34 -69497 50 -69463
rect -50 -69535 50 -69497
rect -50 -70573 50 -70535
rect -50 -70607 -34 -70573
rect 34 -70607 50 -70573
rect -50 -70623 50 -70607
rect -50 -70681 50 -70665
rect -50 -70715 -34 -70681
rect 34 -70715 50 -70681
rect -50 -70753 50 -70715
rect -50 -71791 50 -71753
rect -50 -71825 -34 -71791
rect 34 -71825 50 -71791
rect -50 -71841 50 -71825
rect -50 -71899 50 -71883
rect -50 -71933 -34 -71899
rect 34 -71933 50 -71899
rect -50 -71971 50 -71933
rect -50 -73009 50 -72971
rect -50 -73043 -34 -73009
rect 34 -73043 50 -73009
rect -50 -73059 50 -73043
rect -50 -73117 50 -73101
rect -50 -73151 -34 -73117
rect 34 -73151 50 -73117
rect -50 -73189 50 -73151
rect -50 -74227 50 -74189
rect -50 -74261 -34 -74227
rect 34 -74261 50 -74227
rect -50 -74277 50 -74261
rect -50 -74335 50 -74319
rect -50 -74369 -34 -74335
rect 34 -74369 50 -74335
rect -50 -74407 50 -74369
rect -50 -75445 50 -75407
rect -50 -75479 -34 -75445
rect 34 -75479 50 -75445
rect -50 -75495 50 -75479
rect -50 -75553 50 -75537
rect -50 -75587 -34 -75553
rect 34 -75587 50 -75553
rect -50 -75625 50 -75587
rect -50 -76663 50 -76625
rect -50 -76697 -34 -76663
rect 34 -76697 50 -76663
rect -50 -76713 50 -76697
rect -50 -76771 50 -76755
rect -50 -76805 -34 -76771
rect 34 -76805 50 -76771
rect -50 -76843 50 -76805
rect -50 -77881 50 -77843
rect -50 -77915 -34 -77881
rect 34 -77915 50 -77881
rect -50 -77931 50 -77915
rect -50 -77989 50 -77973
rect -50 -78023 -34 -77989
rect 34 -78023 50 -77989
rect -50 -78061 50 -78023
rect -50 -79099 50 -79061
rect -50 -79133 -34 -79099
rect 34 -79133 50 -79099
rect -50 -79149 50 -79133
rect -50 -79207 50 -79191
rect -50 -79241 -34 -79207
rect 34 -79241 50 -79207
rect -50 -79279 50 -79241
rect -50 -80317 50 -80279
rect -50 -80351 -34 -80317
rect 34 -80351 50 -80317
rect -50 -80367 50 -80351
rect -50 -80425 50 -80409
rect -50 -80459 -34 -80425
rect 34 -80459 50 -80425
rect -50 -80497 50 -80459
rect -50 -81535 50 -81497
rect -50 -81569 -34 -81535
rect 34 -81569 50 -81535
rect -50 -81585 50 -81569
rect -50 -81643 50 -81627
rect -50 -81677 -34 -81643
rect 34 -81677 50 -81643
rect -50 -81715 50 -81677
rect -50 -82753 50 -82715
rect -50 -82787 -34 -82753
rect 34 -82787 50 -82753
rect -50 -82803 50 -82787
rect -50 -82861 50 -82845
rect -50 -82895 -34 -82861
rect 34 -82895 50 -82861
rect -50 -82933 50 -82895
rect -50 -83971 50 -83933
rect -50 -84005 -34 -83971
rect 34 -84005 50 -83971
rect -50 -84021 50 -84005
rect -50 -84079 50 -84063
rect -50 -84113 -34 -84079
rect 34 -84113 50 -84079
rect -50 -84151 50 -84113
rect -50 -85189 50 -85151
rect -50 -85223 -34 -85189
rect 34 -85223 50 -85189
rect -50 -85239 50 -85223
rect -50 -85297 50 -85281
rect -50 -85331 -34 -85297
rect 34 -85331 50 -85297
rect -50 -85369 50 -85331
rect -50 -86407 50 -86369
rect -50 -86441 -34 -86407
rect 34 -86441 50 -86407
rect -50 -86457 50 -86441
rect -50 -86515 50 -86499
rect -50 -86549 -34 -86515
rect 34 -86549 50 -86515
rect -50 -86587 50 -86549
rect -50 -87625 50 -87587
rect -50 -87659 -34 -87625
rect 34 -87659 50 -87625
rect -50 -87675 50 -87659
rect -50 -87733 50 -87717
rect -50 -87767 -34 -87733
rect 34 -87767 50 -87733
rect -50 -87805 50 -87767
rect -50 -88843 50 -88805
rect -50 -88877 -34 -88843
rect 34 -88877 50 -88843
rect -50 -88893 50 -88877
rect -50 -88951 50 -88935
rect -50 -88985 -34 -88951
rect 34 -88985 50 -88951
rect -50 -89023 50 -88985
rect -50 -90061 50 -90023
rect -50 -90095 -34 -90061
rect 34 -90095 50 -90061
rect -50 -90111 50 -90095
rect -50 -90169 50 -90153
rect -50 -90203 -34 -90169
rect 34 -90203 50 -90169
rect -50 -90241 50 -90203
rect -50 -91279 50 -91241
rect -50 -91313 -34 -91279
rect 34 -91313 50 -91279
rect -50 -91329 50 -91313
rect -50 -91387 50 -91371
rect -50 -91421 -34 -91387
rect 34 -91421 50 -91387
rect -50 -91459 50 -91421
rect -50 -92497 50 -92459
rect -50 -92531 -34 -92497
rect 34 -92531 50 -92497
rect -50 -92547 50 -92531
rect -50 -92605 50 -92589
rect -50 -92639 -34 -92605
rect 34 -92639 50 -92605
rect -50 -92677 50 -92639
rect -50 -93715 50 -93677
rect -50 -93749 -34 -93715
rect 34 -93749 50 -93715
rect -50 -93765 50 -93749
rect -50 -93823 50 -93807
rect -50 -93857 -34 -93823
rect 34 -93857 50 -93823
rect -50 -93895 50 -93857
rect -50 -94933 50 -94895
rect -50 -94967 -34 -94933
rect 34 -94967 50 -94933
rect -50 -94983 50 -94967
rect -50 -95041 50 -95025
rect -50 -95075 -34 -95041
rect 34 -95075 50 -95041
rect -50 -95113 50 -95075
rect -50 -96151 50 -96113
rect -50 -96185 -34 -96151
rect 34 -96185 50 -96151
rect -50 -96201 50 -96185
rect -50 -96259 50 -96243
rect -50 -96293 -34 -96259
rect 34 -96293 50 -96259
rect -50 -96331 50 -96293
rect -50 -97369 50 -97331
rect -50 -97403 -34 -97369
rect 34 -97403 50 -97369
rect -50 -97419 50 -97403
rect -50 -97477 50 -97461
rect -50 -97511 -34 -97477
rect 34 -97511 50 -97477
rect -50 -97549 50 -97511
rect -50 -98587 50 -98549
rect -50 -98621 -34 -98587
rect 34 -98621 50 -98587
rect -50 -98637 50 -98621
rect -50 -98695 50 -98679
rect -50 -98729 -34 -98695
rect 34 -98729 50 -98695
rect -50 -98767 50 -98729
rect -50 -99805 50 -99767
rect -50 -99839 -34 -99805
rect 34 -99839 50 -99805
rect -50 -99855 50 -99839
rect -50 -99913 50 -99897
rect -50 -99947 -34 -99913
rect 34 -99947 50 -99913
rect -50 -99985 50 -99947
rect -50 -101023 50 -100985
rect -50 -101057 -34 -101023
rect 34 -101057 50 -101023
rect -50 -101073 50 -101057
rect -50 -101131 50 -101115
rect -50 -101165 -34 -101131
rect 34 -101165 50 -101131
rect -50 -101203 50 -101165
rect -50 -102241 50 -102203
rect -50 -102275 -34 -102241
rect 34 -102275 50 -102241
rect -50 -102291 50 -102275
rect -50 -102349 50 -102333
rect -50 -102383 -34 -102349
rect 34 -102383 50 -102349
rect -50 -102421 50 -102383
rect -50 -103459 50 -103421
rect -50 -103493 -34 -103459
rect 34 -103493 50 -103459
rect -50 -103509 50 -103493
rect -50 -103567 50 -103551
rect -50 -103601 -34 -103567
rect 34 -103601 50 -103567
rect -50 -103639 50 -103601
rect -50 -104677 50 -104639
rect -50 -104711 -34 -104677
rect 34 -104711 50 -104677
rect -50 -104727 50 -104711
rect -50 -104785 50 -104769
rect -50 -104819 -34 -104785
rect 34 -104819 50 -104785
rect -50 -104857 50 -104819
rect -50 -105895 50 -105857
rect -50 -105929 -34 -105895
rect 34 -105929 50 -105895
rect -50 -105945 50 -105929
rect -50 -106003 50 -105987
rect -50 -106037 -34 -106003
rect 34 -106037 50 -106003
rect -50 -106075 50 -106037
rect -50 -107113 50 -107075
rect -50 -107147 -34 -107113
rect 34 -107147 50 -107113
rect -50 -107163 50 -107147
rect -50 -107221 50 -107205
rect -50 -107255 -34 -107221
rect 34 -107255 50 -107221
rect -50 -107293 50 -107255
rect -50 -108331 50 -108293
rect -50 -108365 -34 -108331
rect 34 -108365 50 -108331
rect -50 -108381 50 -108365
rect -50 -108439 50 -108423
rect -50 -108473 -34 -108439
rect 34 -108473 50 -108439
rect -50 -108511 50 -108473
rect -50 -109549 50 -109511
rect -50 -109583 -34 -109549
rect 34 -109583 50 -109549
rect -50 -109599 50 -109583
rect -50 -109657 50 -109641
rect -50 -109691 -34 -109657
rect 34 -109691 50 -109657
rect -50 -109729 50 -109691
rect -50 -110767 50 -110729
rect -50 -110801 -34 -110767
rect 34 -110801 50 -110767
rect -50 -110817 50 -110801
rect -50 -110875 50 -110859
rect -50 -110909 -34 -110875
rect 34 -110909 50 -110875
rect -50 -110947 50 -110909
rect -50 -111985 50 -111947
rect -50 -112019 -34 -111985
rect 34 -112019 50 -111985
rect -50 -112035 50 -112019
rect -50 -112093 50 -112077
rect -50 -112127 -34 -112093
rect 34 -112127 50 -112093
rect -50 -112165 50 -112127
rect -50 -113203 50 -113165
rect -50 -113237 -34 -113203
rect 34 -113237 50 -113203
rect -50 -113253 50 -113237
rect -50 -113311 50 -113295
rect -50 -113345 -34 -113311
rect 34 -113345 50 -113311
rect -50 -113383 50 -113345
rect -50 -114421 50 -114383
rect -50 -114455 -34 -114421
rect 34 -114455 50 -114421
rect -50 -114471 50 -114455
rect -50 -114529 50 -114513
rect -50 -114563 -34 -114529
rect 34 -114563 50 -114529
rect -50 -114601 50 -114563
rect -50 -115639 50 -115601
rect -50 -115673 -34 -115639
rect 34 -115673 50 -115639
rect -50 -115689 50 -115673
rect -50 -115747 50 -115731
rect -50 -115781 -34 -115747
rect 34 -115781 50 -115747
rect -50 -115819 50 -115781
rect -50 -116857 50 -116819
rect -50 -116891 -34 -116857
rect 34 -116891 50 -116857
rect -50 -116907 50 -116891
rect -50 -116965 50 -116949
rect -50 -116999 -34 -116965
rect 34 -116999 50 -116965
rect -50 -117037 50 -116999
rect -50 -118075 50 -118037
rect -50 -118109 -34 -118075
rect 34 -118109 50 -118075
rect -50 -118125 50 -118109
rect -50 -118183 50 -118167
rect -50 -118217 -34 -118183
rect 34 -118217 50 -118183
rect -50 -118255 50 -118217
rect -50 -119293 50 -119255
rect -50 -119327 -34 -119293
rect 34 -119327 50 -119293
rect -50 -119343 50 -119327
rect -50 -119401 50 -119385
rect -50 -119435 -34 -119401
rect 34 -119435 50 -119401
rect -50 -119473 50 -119435
rect -50 -120511 50 -120473
rect -50 -120545 -34 -120511
rect 34 -120545 50 -120511
rect -50 -120561 50 -120545
rect -50 -120619 50 -120603
rect -50 -120653 -34 -120619
rect 34 -120653 50 -120619
rect -50 -120691 50 -120653
rect -50 -121729 50 -121691
rect -50 -121763 -34 -121729
rect 34 -121763 50 -121729
rect -50 -121779 50 -121763
rect -50 -121837 50 -121821
rect -50 -121871 -34 -121837
rect 34 -121871 50 -121837
rect -50 -121909 50 -121871
rect -50 -122947 50 -122909
rect -50 -122981 -34 -122947
rect 34 -122981 50 -122947
rect -50 -122997 50 -122981
rect -50 -123055 50 -123039
rect -50 -123089 -34 -123055
rect 34 -123089 50 -123055
rect -50 -123127 50 -123089
rect -50 -124165 50 -124127
rect -50 -124199 -34 -124165
rect 34 -124199 50 -124165
rect -50 -124215 50 -124199
rect -50 -124273 50 -124257
rect -50 -124307 -34 -124273
rect 34 -124307 50 -124273
rect -50 -124345 50 -124307
rect -50 -125383 50 -125345
rect -50 -125417 -34 -125383
rect 34 -125417 50 -125383
rect -50 -125433 50 -125417
rect -50 -125491 50 -125475
rect -50 -125525 -34 -125491
rect 34 -125525 50 -125491
rect -50 -125563 50 -125525
rect -50 -126601 50 -126563
rect -50 -126635 -34 -126601
rect 34 -126635 50 -126601
rect -50 -126651 50 -126635
rect -50 -126709 50 -126693
rect -50 -126743 -34 -126709
rect 34 -126743 50 -126709
rect -50 -126781 50 -126743
rect -50 -127819 50 -127781
rect -50 -127853 -34 -127819
rect 34 -127853 50 -127819
rect -50 -127869 50 -127853
rect -50 -127927 50 -127911
rect -50 -127961 -34 -127927
rect 34 -127961 50 -127927
rect -50 -127999 50 -127961
rect -50 -129037 50 -128999
rect -50 -129071 -34 -129037
rect 34 -129071 50 -129037
rect -50 -129087 50 -129071
rect -50 -129145 50 -129129
rect -50 -129179 -34 -129145
rect 34 -129179 50 -129145
rect -50 -129217 50 -129179
rect -50 -130255 50 -130217
rect -50 -130289 -34 -130255
rect 34 -130289 50 -130255
rect -50 -130305 50 -130289
rect -50 -130363 50 -130347
rect -50 -130397 -34 -130363
rect 34 -130397 50 -130363
rect -50 -130435 50 -130397
rect -50 -131473 50 -131435
rect -50 -131507 -34 -131473
rect 34 -131507 50 -131473
rect -50 -131523 50 -131507
rect -50 -131581 50 -131565
rect -50 -131615 -34 -131581
rect 34 -131615 50 -131581
rect -50 -131653 50 -131615
rect -50 -132691 50 -132653
rect -50 -132725 -34 -132691
rect 34 -132725 50 -132691
rect -50 -132741 50 -132725
rect -50 -132799 50 -132783
rect -50 -132833 -34 -132799
rect 34 -132833 50 -132799
rect -50 -132871 50 -132833
rect -50 -133909 50 -133871
rect -50 -133943 -34 -133909
rect 34 -133943 50 -133909
rect -50 -133959 50 -133943
rect -50 -134017 50 -134001
rect -50 -134051 -34 -134017
rect 34 -134051 50 -134017
rect -50 -134089 50 -134051
rect -50 -135127 50 -135089
rect -50 -135161 -34 -135127
rect 34 -135161 50 -135127
rect -50 -135177 50 -135161
rect -50 -135235 50 -135219
rect -50 -135269 -34 -135235
rect 34 -135269 50 -135235
rect -50 -135307 50 -135269
rect -50 -136345 50 -136307
rect -50 -136379 -34 -136345
rect 34 -136379 50 -136345
rect -50 -136395 50 -136379
rect -50 -136453 50 -136437
rect -50 -136487 -34 -136453
rect 34 -136487 50 -136453
rect -50 -136525 50 -136487
rect -50 -137563 50 -137525
rect -50 -137597 -34 -137563
rect 34 -137597 50 -137563
rect -50 -137613 50 -137597
rect -50 -137671 50 -137655
rect -50 -137705 -34 -137671
rect 34 -137705 50 -137671
rect -50 -137743 50 -137705
rect -50 -138781 50 -138743
rect -50 -138815 -34 -138781
rect 34 -138815 50 -138781
rect -50 -138831 50 -138815
rect -50 -138889 50 -138873
rect -50 -138923 -34 -138889
rect 34 -138923 50 -138889
rect -50 -138961 50 -138923
rect -50 -139999 50 -139961
rect -50 -140033 -34 -139999
rect 34 -140033 50 -139999
rect -50 -140049 50 -140033
rect -50 -140107 50 -140091
rect -50 -140141 -34 -140107
rect 34 -140141 50 -140107
rect -50 -140179 50 -140141
rect -50 -141217 50 -141179
rect -50 -141251 -34 -141217
rect 34 -141251 50 -141217
rect -50 -141267 50 -141251
rect -50 -141325 50 -141309
rect -50 -141359 -34 -141325
rect 34 -141359 50 -141325
rect -50 -141397 50 -141359
rect -50 -142435 50 -142397
rect -50 -142469 -34 -142435
rect 34 -142469 50 -142435
rect -50 -142485 50 -142469
rect -50 -142543 50 -142527
rect -50 -142577 -34 -142543
rect 34 -142577 50 -142543
rect -50 -142615 50 -142577
rect -50 -143653 50 -143615
rect -50 -143687 -34 -143653
rect 34 -143687 50 -143653
rect -50 -143703 50 -143687
rect -50 -143761 50 -143745
rect -50 -143795 -34 -143761
rect 34 -143795 50 -143761
rect -50 -143833 50 -143795
rect -50 -144871 50 -144833
rect -50 -144905 -34 -144871
rect 34 -144905 50 -144871
rect -50 -144921 50 -144905
rect -50 -144979 50 -144963
rect -50 -145013 -34 -144979
rect 34 -145013 50 -144979
rect -50 -145051 50 -145013
rect -50 -146089 50 -146051
rect -50 -146123 -34 -146089
rect 34 -146123 50 -146089
rect -50 -146139 50 -146123
rect -50 -146197 50 -146181
rect -50 -146231 -34 -146197
rect 34 -146231 50 -146197
rect -50 -146269 50 -146231
rect -50 -147307 50 -147269
rect -50 -147341 -34 -147307
rect 34 -147341 50 -147307
rect -50 -147357 50 -147341
rect -50 -147415 50 -147399
rect -50 -147449 -34 -147415
rect 34 -147449 50 -147415
rect -50 -147487 50 -147449
rect -50 -148525 50 -148487
rect -50 -148559 -34 -148525
rect 34 -148559 50 -148525
rect -50 -148575 50 -148559
rect -50 -148633 50 -148617
rect -50 -148667 -34 -148633
rect 34 -148667 50 -148633
rect -50 -148705 50 -148667
rect -50 -149743 50 -149705
rect -50 -149777 -34 -149743
rect 34 -149777 50 -149743
rect -50 -149793 50 -149777
rect -50 -149851 50 -149835
rect -50 -149885 -34 -149851
rect 34 -149885 50 -149851
rect -50 -149923 50 -149885
rect -50 -150961 50 -150923
rect -50 -150995 -34 -150961
rect 34 -150995 50 -150961
rect -50 -151011 50 -150995
rect -50 -151069 50 -151053
rect -50 -151103 -34 -151069
rect 34 -151103 50 -151069
rect -50 -151141 50 -151103
rect -50 -152179 50 -152141
rect -50 -152213 -34 -152179
rect 34 -152213 50 -152179
rect -50 -152229 50 -152213
rect -50 -152287 50 -152271
rect -50 -152321 -34 -152287
rect 34 -152321 50 -152287
rect -50 -152359 50 -152321
rect -50 -153397 50 -153359
rect -50 -153431 -34 -153397
rect 34 -153431 50 -153397
rect -50 -153447 50 -153431
rect -50 -153505 50 -153489
rect -50 -153539 -34 -153505
rect 34 -153539 50 -153505
rect -50 -153577 50 -153539
rect -50 -154615 50 -154577
rect -50 -154649 -34 -154615
rect 34 -154649 50 -154615
rect -50 -154665 50 -154649
rect -50 -154723 50 -154707
rect -50 -154757 -34 -154723
rect 34 -154757 50 -154723
rect -50 -154795 50 -154757
rect -50 -155833 50 -155795
rect -50 -155867 -34 -155833
rect 34 -155867 50 -155833
rect -50 -155883 50 -155867
rect -50 -155941 50 -155925
rect -50 -155975 -34 -155941
rect 34 -155975 50 -155941
rect -50 -156013 50 -155975
rect -50 -157051 50 -157013
rect -50 -157085 -34 -157051
rect 34 -157085 50 -157051
rect -50 -157101 50 -157085
rect -50 -157159 50 -157143
rect -50 -157193 -34 -157159
rect 34 -157193 50 -157159
rect -50 -157231 50 -157193
rect -50 -158269 50 -158231
rect -50 -158303 -34 -158269
rect 34 -158303 50 -158269
rect -50 -158319 50 -158303
rect -50 -158377 50 -158361
rect -50 -158411 -34 -158377
rect 34 -158411 50 -158377
rect -50 -158449 50 -158411
rect -50 -159487 50 -159449
rect -50 -159521 -34 -159487
rect 34 -159521 50 -159487
rect -50 -159537 50 -159521
rect -50 -159595 50 -159579
rect -50 -159629 -34 -159595
rect 34 -159629 50 -159595
rect -50 -159667 50 -159629
rect -50 -160705 50 -160667
rect -50 -160739 -34 -160705
rect 34 -160739 50 -160705
rect -50 -160755 50 -160739
rect -50 -160813 50 -160797
rect -50 -160847 -34 -160813
rect 34 -160847 50 -160813
rect -50 -160885 50 -160847
rect -50 -161923 50 -161885
rect -50 -161957 -34 -161923
rect 34 -161957 50 -161923
rect -50 -161973 50 -161957
rect -50 -162031 50 -162015
rect -50 -162065 -34 -162031
rect 34 -162065 50 -162031
rect -50 -162103 50 -162065
rect -50 -163141 50 -163103
rect -50 -163175 -34 -163141
rect 34 -163175 50 -163141
rect -50 -163191 50 -163175
rect -50 -163249 50 -163233
rect -50 -163283 -34 -163249
rect 34 -163283 50 -163249
rect -50 -163321 50 -163283
rect -50 -164359 50 -164321
rect -50 -164393 -34 -164359
rect 34 -164393 50 -164359
rect -50 -164409 50 -164393
rect -50 -164467 50 -164451
rect -50 -164501 -34 -164467
rect 34 -164501 50 -164467
rect -50 -164539 50 -164501
rect -50 -165577 50 -165539
rect -50 -165611 -34 -165577
rect 34 -165611 50 -165577
rect -50 -165627 50 -165611
rect -50 -165685 50 -165669
rect -50 -165719 -34 -165685
rect 34 -165719 50 -165685
rect -50 -165757 50 -165719
rect -50 -166795 50 -166757
rect -50 -166829 -34 -166795
rect 34 -166829 50 -166795
rect -50 -166845 50 -166829
rect -50 -166903 50 -166887
rect -50 -166937 -34 -166903
rect 34 -166937 50 -166903
rect -50 -166975 50 -166937
rect -50 -168013 50 -167975
rect -50 -168047 -34 -168013
rect 34 -168047 50 -168013
rect -50 -168063 50 -168047
rect -50 -168121 50 -168105
rect -50 -168155 -34 -168121
rect 34 -168155 50 -168121
rect -50 -168193 50 -168155
rect -50 -169231 50 -169193
rect -50 -169265 -34 -169231
rect 34 -169265 50 -169231
rect -50 -169281 50 -169265
rect -50 -169339 50 -169323
rect -50 -169373 -34 -169339
rect 34 -169373 50 -169339
rect -50 -169411 50 -169373
rect -50 -170449 50 -170411
rect -50 -170483 -34 -170449
rect 34 -170483 50 -170449
rect -50 -170499 50 -170483
rect -50 -170557 50 -170541
rect -50 -170591 -34 -170557
rect 34 -170591 50 -170557
rect -50 -170629 50 -170591
rect -50 -171667 50 -171629
rect -50 -171701 -34 -171667
rect 34 -171701 50 -171667
rect -50 -171717 50 -171701
rect -50 -171775 50 -171759
rect -50 -171809 -34 -171775
rect 34 -171809 50 -171775
rect -50 -171847 50 -171809
rect -50 -172885 50 -172847
rect -50 -172919 -34 -172885
rect 34 -172919 50 -172885
rect -50 -172935 50 -172919
rect -50 -172993 50 -172977
rect -50 -173027 -34 -172993
rect 34 -173027 50 -172993
rect -50 -173065 50 -173027
rect -50 -174103 50 -174065
rect -50 -174137 -34 -174103
rect 34 -174137 50 -174103
rect -50 -174153 50 -174137
rect -50 -174211 50 -174195
rect -50 -174245 -34 -174211
rect 34 -174245 50 -174211
rect -50 -174283 50 -174245
rect -50 -175321 50 -175283
rect -50 -175355 -34 -175321
rect 34 -175355 50 -175321
rect -50 -175371 50 -175355
rect -50 -175429 50 -175413
rect -50 -175463 -34 -175429
rect 34 -175463 50 -175429
rect -50 -175501 50 -175463
rect -50 -176539 50 -176501
rect -50 -176573 -34 -176539
rect 34 -176573 50 -176539
rect -50 -176589 50 -176573
rect -50 -176647 50 -176631
rect -50 -176681 -34 -176647
rect 34 -176681 50 -176647
rect -50 -176719 50 -176681
rect -50 -177757 50 -177719
rect -50 -177791 -34 -177757
rect 34 -177791 50 -177757
rect -50 -177807 50 -177791
rect -50 -177865 50 -177849
rect -50 -177899 -34 -177865
rect 34 -177899 50 -177865
rect -50 -177937 50 -177899
rect -50 -178975 50 -178937
rect -50 -179009 -34 -178975
rect 34 -179009 50 -178975
rect -50 -179025 50 -179009
rect -50 -179083 50 -179067
rect -50 -179117 -34 -179083
rect 34 -179117 50 -179083
rect -50 -179155 50 -179117
rect -50 -180193 50 -180155
rect -50 -180227 -34 -180193
rect 34 -180227 50 -180193
rect -50 -180243 50 -180227
rect -50 -180301 50 -180285
rect -50 -180335 -34 -180301
rect 34 -180335 50 -180301
rect -50 -180373 50 -180335
rect -50 -181411 50 -181373
rect -50 -181445 -34 -181411
rect 34 -181445 50 -181411
rect -50 -181461 50 -181445
rect -50 -181519 50 -181503
rect -50 -181553 -34 -181519
rect 34 -181553 50 -181519
rect -50 -181591 50 -181553
rect -50 -182629 50 -182591
rect -50 -182663 -34 -182629
rect 34 -182663 50 -182629
rect -50 -182679 50 -182663
rect -50 -182737 50 -182721
rect -50 -182771 -34 -182737
rect 34 -182771 50 -182737
rect -50 -182809 50 -182771
rect -50 -183847 50 -183809
rect -50 -183881 -34 -183847
rect 34 -183881 50 -183847
rect -50 -183897 50 -183881
rect -50 -183955 50 -183939
rect -50 -183989 -34 -183955
rect 34 -183989 50 -183955
rect -50 -184027 50 -183989
rect -50 -185065 50 -185027
rect -50 -185099 -34 -185065
rect 34 -185099 50 -185065
rect -50 -185115 50 -185099
rect -50 -185173 50 -185157
rect -50 -185207 -34 -185173
rect 34 -185207 50 -185173
rect -50 -185245 50 -185207
rect -50 -186283 50 -186245
rect -50 -186317 -34 -186283
rect 34 -186317 50 -186283
rect -50 -186333 50 -186317
rect -50 -186391 50 -186375
rect -50 -186425 -34 -186391
rect 34 -186425 50 -186391
rect -50 -186463 50 -186425
rect -50 -187501 50 -187463
rect -50 -187535 -34 -187501
rect 34 -187535 50 -187501
rect -50 -187551 50 -187535
rect -50 -187609 50 -187593
rect -50 -187643 -34 -187609
rect 34 -187643 50 -187609
rect -50 -187681 50 -187643
rect -50 -188719 50 -188681
rect -50 -188753 -34 -188719
rect 34 -188753 50 -188719
rect -50 -188769 50 -188753
rect -50 -188827 50 -188811
rect -50 -188861 -34 -188827
rect 34 -188861 50 -188827
rect -50 -188899 50 -188861
rect -50 -189937 50 -189899
rect -50 -189971 -34 -189937
rect 34 -189971 50 -189937
rect -50 -189987 50 -189971
rect -50 -190045 50 -190029
rect -50 -190079 -34 -190045
rect 34 -190079 50 -190045
rect -50 -190117 50 -190079
rect -50 -191155 50 -191117
rect -50 -191189 -34 -191155
rect 34 -191189 50 -191155
rect -50 -191205 50 -191189
rect -50 -191263 50 -191247
rect -50 -191297 -34 -191263
rect 34 -191297 50 -191263
rect -50 -191335 50 -191297
rect -50 -192373 50 -192335
rect -50 -192407 -34 -192373
rect 34 -192407 50 -192373
rect -50 -192423 50 -192407
rect -50 -192481 50 -192465
rect -50 -192515 -34 -192481
rect 34 -192515 50 -192481
rect -50 -192553 50 -192515
rect -50 -193591 50 -193553
rect -50 -193625 -34 -193591
rect 34 -193625 50 -193591
rect -50 -193641 50 -193625
rect -50 -193699 50 -193683
rect -50 -193733 -34 -193699
rect 34 -193733 50 -193699
rect -50 -193771 50 -193733
rect -50 -194809 50 -194771
rect -50 -194843 -34 -194809
rect 34 -194843 50 -194809
rect -50 -194859 50 -194843
rect -50 -194917 50 -194901
rect -50 -194951 -34 -194917
rect 34 -194951 50 -194917
rect -50 -194989 50 -194951
rect -50 -196027 50 -195989
rect -50 -196061 -34 -196027
rect 34 -196061 50 -196027
rect -50 -196077 50 -196061
rect -50 -196135 50 -196119
rect -50 -196169 -34 -196135
rect 34 -196169 50 -196135
rect -50 -196207 50 -196169
rect -50 -197245 50 -197207
rect -50 -197279 -34 -197245
rect 34 -197279 50 -197245
rect -50 -197295 50 -197279
rect -50 -197353 50 -197337
rect -50 -197387 -34 -197353
rect 34 -197387 50 -197353
rect -50 -197425 50 -197387
rect -50 -198463 50 -198425
rect -50 -198497 -34 -198463
rect 34 -198497 50 -198463
rect -50 -198513 50 -198497
rect -50 -198571 50 -198555
rect -50 -198605 -34 -198571
rect 34 -198605 50 -198571
rect -50 -198643 50 -198605
rect -50 -199681 50 -199643
rect -50 -199715 -34 -199681
rect 34 -199715 50 -199681
rect -50 -199731 50 -199715
rect -50 -199789 50 -199773
rect -50 -199823 -34 -199789
rect 34 -199823 50 -199789
rect -50 -199861 50 -199823
rect -50 -200899 50 -200861
rect -50 -200933 -34 -200899
rect 34 -200933 50 -200899
rect -50 -200949 50 -200933
rect -50 -201007 50 -200991
rect -50 -201041 -34 -201007
rect 34 -201041 50 -201007
rect -50 -201079 50 -201041
rect -50 -202117 50 -202079
rect -50 -202151 -34 -202117
rect 34 -202151 50 -202117
rect -50 -202167 50 -202151
rect -50 -202225 50 -202209
rect -50 -202259 -34 -202225
rect 34 -202259 50 -202225
rect -50 -202297 50 -202259
rect -50 -203335 50 -203297
rect -50 -203369 -34 -203335
rect 34 -203369 50 -203335
rect -50 -203385 50 -203369
rect -50 -203443 50 -203427
rect -50 -203477 -34 -203443
rect 34 -203477 50 -203443
rect -50 -203515 50 -203477
rect -50 -204553 50 -204515
rect -50 -204587 -34 -204553
rect 34 -204587 50 -204553
rect -50 -204603 50 -204587
rect -50 -204661 50 -204645
rect -50 -204695 -34 -204661
rect 34 -204695 50 -204661
rect -50 -204733 50 -204695
rect -50 -205771 50 -205733
rect -50 -205805 -34 -205771
rect 34 -205805 50 -205771
rect -50 -205821 50 -205805
rect -50 -205879 50 -205863
rect -50 -205913 -34 -205879
rect 34 -205913 50 -205879
rect -50 -205951 50 -205913
rect -50 -206989 50 -206951
rect -50 -207023 -34 -206989
rect 34 -207023 50 -206989
rect -50 -207039 50 -207023
rect -50 -207097 50 -207081
rect -50 -207131 -34 -207097
rect 34 -207131 50 -207097
rect -50 -207169 50 -207131
rect -50 -208207 50 -208169
rect -50 -208241 -34 -208207
rect 34 -208241 50 -208207
rect -50 -208257 50 -208241
rect -50 -208315 50 -208299
rect -50 -208349 -34 -208315
rect 34 -208349 50 -208315
rect -50 -208387 50 -208349
rect -50 -209425 50 -209387
rect -50 -209459 -34 -209425
rect 34 -209459 50 -209425
rect -50 -209475 50 -209459
rect -50 -209533 50 -209517
rect -50 -209567 -34 -209533
rect 34 -209567 50 -209533
rect -50 -209605 50 -209567
rect -50 -210643 50 -210605
rect -50 -210677 -34 -210643
rect 34 -210677 50 -210643
rect -50 -210693 50 -210677
rect -50 -210751 50 -210735
rect -50 -210785 -34 -210751
rect 34 -210785 50 -210751
rect -50 -210823 50 -210785
rect -50 -211861 50 -211823
rect -50 -211895 -34 -211861
rect 34 -211895 50 -211861
rect -50 -211911 50 -211895
rect -50 -211969 50 -211953
rect -50 -212003 -34 -211969
rect 34 -212003 50 -211969
rect -50 -212041 50 -212003
rect -50 -213079 50 -213041
rect -50 -213113 -34 -213079
rect 34 -213113 50 -213079
rect -50 -213129 50 -213113
rect -50 -213187 50 -213171
rect -50 -213221 -34 -213187
rect 34 -213221 50 -213187
rect -50 -213259 50 -213221
rect -50 -214297 50 -214259
rect -50 -214331 -34 -214297
rect 34 -214331 50 -214297
rect -50 -214347 50 -214331
rect -50 -214405 50 -214389
rect -50 -214439 -34 -214405
rect 34 -214439 50 -214405
rect -50 -214477 50 -214439
rect -50 -215515 50 -215477
rect -50 -215549 -34 -215515
rect 34 -215549 50 -215515
rect -50 -215565 50 -215549
rect -50 -215623 50 -215607
rect -50 -215657 -34 -215623
rect 34 -215657 50 -215623
rect -50 -215695 50 -215657
rect -50 -216733 50 -216695
rect -50 -216767 -34 -216733
rect 34 -216767 50 -216733
rect -50 -216783 50 -216767
rect -50 -216841 50 -216825
rect -50 -216875 -34 -216841
rect 34 -216875 50 -216841
rect -50 -216913 50 -216875
rect -50 -217951 50 -217913
rect -50 -217985 -34 -217951
rect 34 -217985 50 -217951
rect -50 -218001 50 -217985
rect -50 -218059 50 -218043
rect -50 -218093 -34 -218059
rect 34 -218093 50 -218059
rect -50 -218131 50 -218093
rect -50 -219169 50 -219131
rect -50 -219203 -34 -219169
rect 34 -219203 50 -219169
rect -50 -219219 50 -219203
rect -50 -219277 50 -219261
rect -50 -219311 -34 -219277
rect 34 -219311 50 -219277
rect -50 -219349 50 -219311
rect -50 -220387 50 -220349
rect -50 -220421 -34 -220387
rect 34 -220421 50 -220387
rect -50 -220437 50 -220421
rect -50 -220495 50 -220479
rect -50 -220529 -34 -220495
rect 34 -220529 50 -220495
rect -50 -220567 50 -220529
rect -50 -221605 50 -221567
rect -50 -221639 -34 -221605
rect 34 -221639 50 -221605
rect -50 -221655 50 -221639
rect -50 -221713 50 -221697
rect -50 -221747 -34 -221713
rect 34 -221747 50 -221713
rect -50 -221785 50 -221747
rect -50 -222823 50 -222785
rect -50 -222857 -34 -222823
rect 34 -222857 50 -222823
rect -50 -222873 50 -222857
rect -50 -222931 50 -222915
rect -50 -222965 -34 -222931
rect 34 -222965 50 -222931
rect -50 -223003 50 -222965
rect -50 -224041 50 -224003
rect -50 -224075 -34 -224041
rect 34 -224075 50 -224041
rect -50 -224091 50 -224075
rect -50 -224149 50 -224133
rect -50 -224183 -34 -224149
rect 34 -224183 50 -224149
rect -50 -224221 50 -224183
rect -50 -225259 50 -225221
rect -50 -225293 -34 -225259
rect 34 -225293 50 -225259
rect -50 -225309 50 -225293
rect -50 -225367 50 -225351
rect -50 -225401 -34 -225367
rect 34 -225401 50 -225367
rect -50 -225439 50 -225401
rect -50 -226477 50 -226439
rect -50 -226511 -34 -226477
rect 34 -226511 50 -226477
rect -50 -226527 50 -226511
rect -50 -226585 50 -226569
rect -50 -226619 -34 -226585
rect 34 -226619 50 -226585
rect -50 -226657 50 -226619
rect -50 -227695 50 -227657
rect -50 -227729 -34 -227695
rect 34 -227729 50 -227695
rect -50 -227745 50 -227729
rect -50 -227803 50 -227787
rect -50 -227837 -34 -227803
rect 34 -227837 50 -227803
rect -50 -227875 50 -227837
rect -50 -228913 50 -228875
rect -50 -228947 -34 -228913
rect 34 -228947 50 -228913
rect -50 -228963 50 -228947
rect -50 -229021 50 -229005
rect -50 -229055 -34 -229021
rect 34 -229055 50 -229021
rect -50 -229093 50 -229055
rect -50 -230131 50 -230093
rect -50 -230165 -34 -230131
rect 34 -230165 50 -230131
rect -50 -230181 50 -230165
rect -50 -230239 50 -230223
rect -50 -230273 -34 -230239
rect 34 -230273 50 -230239
rect -50 -230311 50 -230273
rect -50 -231349 50 -231311
rect -50 -231383 -34 -231349
rect 34 -231383 50 -231349
rect -50 -231399 50 -231383
rect -50 -231457 50 -231441
rect -50 -231491 -34 -231457
rect 34 -231491 50 -231457
rect -50 -231529 50 -231491
rect -50 -232567 50 -232529
rect -50 -232601 -34 -232567
rect 34 -232601 50 -232567
rect -50 -232617 50 -232601
rect -50 -232675 50 -232659
rect -50 -232709 -34 -232675
rect 34 -232709 50 -232675
rect -50 -232747 50 -232709
rect -50 -233785 50 -233747
rect -50 -233819 -34 -233785
rect 34 -233819 50 -233785
rect -50 -233835 50 -233819
rect -50 -233893 50 -233877
rect -50 -233927 -34 -233893
rect 34 -233927 50 -233893
rect -50 -233965 50 -233927
rect -50 -235003 50 -234965
rect -50 -235037 -34 -235003
rect 34 -235037 50 -235003
rect -50 -235053 50 -235037
rect -50 -235111 50 -235095
rect -50 -235145 -34 -235111
rect 34 -235145 50 -235111
rect -50 -235183 50 -235145
rect -50 -236221 50 -236183
rect -50 -236255 -34 -236221
rect 34 -236255 50 -236221
rect -50 -236271 50 -236255
rect -50 -236329 50 -236313
rect -50 -236363 -34 -236329
rect 34 -236363 50 -236329
rect -50 -236401 50 -236363
rect -50 -237439 50 -237401
rect -50 -237473 -34 -237439
rect 34 -237473 50 -237439
rect -50 -237489 50 -237473
rect -50 -237547 50 -237531
rect -50 -237581 -34 -237547
rect 34 -237581 50 -237547
rect -50 -237619 50 -237581
rect -50 -238657 50 -238619
rect -50 -238691 -34 -238657
rect 34 -238691 50 -238657
rect -50 -238707 50 -238691
rect -50 -238765 50 -238749
rect -50 -238799 -34 -238765
rect 34 -238799 50 -238765
rect -50 -238837 50 -238799
rect -50 -239875 50 -239837
rect -50 -239909 -34 -239875
rect 34 -239909 50 -239875
rect -50 -239925 50 -239909
rect -50 -239983 50 -239967
rect -50 -240017 -34 -239983
rect 34 -240017 50 -239983
rect -50 -240055 50 -240017
rect -50 -241093 50 -241055
rect -50 -241127 -34 -241093
rect 34 -241127 50 -241093
rect -50 -241143 50 -241127
rect -50 -241201 50 -241185
rect -50 -241235 -34 -241201
rect 34 -241235 50 -241201
rect -50 -241273 50 -241235
rect -50 -242311 50 -242273
rect -50 -242345 -34 -242311
rect 34 -242345 50 -242311
rect -50 -242361 50 -242345
rect -50 -242419 50 -242403
rect -50 -242453 -34 -242419
rect 34 -242453 50 -242419
rect -50 -242491 50 -242453
rect -50 -243529 50 -243491
rect -50 -243563 -34 -243529
rect 34 -243563 50 -243529
rect -50 -243579 50 -243563
rect -50 -243637 50 -243621
rect -50 -243671 -34 -243637
rect 34 -243671 50 -243637
rect -50 -243709 50 -243671
rect -50 -244747 50 -244709
rect -50 -244781 -34 -244747
rect 34 -244781 50 -244747
rect -50 -244797 50 -244781
rect -50 -244855 50 -244839
rect -50 -244889 -34 -244855
rect 34 -244889 50 -244855
rect -50 -244927 50 -244889
rect -50 -245965 50 -245927
rect -50 -245999 -34 -245965
rect 34 -245999 50 -245965
rect -50 -246015 50 -245999
rect -50 -246073 50 -246057
rect -50 -246107 -34 -246073
rect 34 -246107 50 -246073
rect -50 -246145 50 -246107
rect -50 -247183 50 -247145
rect -50 -247217 -34 -247183
rect 34 -247217 50 -247183
rect -50 -247233 50 -247217
rect -50 -247291 50 -247275
rect -50 -247325 -34 -247291
rect 34 -247325 50 -247291
rect -50 -247363 50 -247325
rect -50 -248401 50 -248363
rect -50 -248435 -34 -248401
rect 34 -248435 50 -248401
rect -50 -248451 50 -248435
rect -50 -248509 50 -248493
rect -50 -248543 -34 -248509
rect 34 -248543 50 -248509
rect -50 -248581 50 -248543
rect -50 -249619 50 -249581
rect -50 -249653 -34 -249619
rect 34 -249653 50 -249619
rect -50 -249669 50 -249653
rect -50 -249727 50 -249711
rect -50 -249761 -34 -249727
rect 34 -249761 50 -249727
rect -50 -249799 50 -249761
rect -50 -250837 50 -250799
rect -50 -250871 -34 -250837
rect 34 -250871 50 -250837
rect -50 -250887 50 -250871
rect -50 -250945 50 -250929
rect -50 -250979 -34 -250945
rect 34 -250979 50 -250945
rect -50 -251017 50 -250979
rect -50 -252055 50 -252017
rect -50 -252089 -34 -252055
rect 34 -252089 50 -252055
rect -50 -252105 50 -252089
rect -50 -252163 50 -252147
rect -50 -252197 -34 -252163
rect 34 -252197 50 -252163
rect -50 -252235 50 -252197
rect -50 -253273 50 -253235
rect -50 -253307 -34 -253273
rect 34 -253307 50 -253273
rect -50 -253323 50 -253307
rect -50 -253381 50 -253365
rect -50 -253415 -34 -253381
rect 34 -253415 50 -253381
rect -50 -253453 50 -253415
rect -50 -254491 50 -254453
rect -50 -254525 -34 -254491
rect 34 -254525 50 -254491
rect -50 -254541 50 -254525
rect -50 -254599 50 -254583
rect -50 -254633 -34 -254599
rect 34 -254633 50 -254599
rect -50 -254671 50 -254633
rect -50 -255709 50 -255671
rect -50 -255743 -34 -255709
rect 34 -255743 50 -255709
rect -50 -255759 50 -255743
rect -50 -255817 50 -255801
rect -50 -255851 -34 -255817
rect 34 -255851 50 -255817
rect -50 -255889 50 -255851
rect -50 -256927 50 -256889
rect -50 -256961 -34 -256927
rect 34 -256961 50 -256927
rect -50 -256977 50 -256961
rect -50 -257035 50 -257019
rect -50 -257069 -34 -257035
rect 34 -257069 50 -257035
rect -50 -257107 50 -257069
rect -50 -258145 50 -258107
rect -50 -258179 -34 -258145
rect 34 -258179 50 -258145
rect -50 -258195 50 -258179
rect -50 -258253 50 -258237
rect -50 -258287 -34 -258253
rect 34 -258287 50 -258253
rect -50 -258325 50 -258287
rect -50 -259363 50 -259325
rect -50 -259397 -34 -259363
rect 34 -259397 50 -259363
rect -50 -259413 50 -259397
rect -50 -259471 50 -259455
rect -50 -259505 -34 -259471
rect 34 -259505 50 -259471
rect -50 -259543 50 -259505
rect -50 -260581 50 -260543
rect -50 -260615 -34 -260581
rect 34 -260615 50 -260581
rect -50 -260631 50 -260615
rect -50 -260689 50 -260673
rect -50 -260723 -34 -260689
rect 34 -260723 50 -260689
rect -50 -260761 50 -260723
rect -50 -261799 50 -261761
rect -50 -261833 -34 -261799
rect 34 -261833 50 -261799
rect -50 -261849 50 -261833
rect -50 -261907 50 -261891
rect -50 -261941 -34 -261907
rect 34 -261941 50 -261907
rect -50 -261979 50 -261941
rect -50 -263017 50 -262979
rect -50 -263051 -34 -263017
rect 34 -263051 50 -263017
rect -50 -263067 50 -263051
rect -50 -263125 50 -263109
rect -50 -263159 -34 -263125
rect 34 -263159 50 -263125
rect -50 -263197 50 -263159
rect -50 -264235 50 -264197
rect -50 -264269 -34 -264235
rect 34 -264269 50 -264235
rect -50 -264285 50 -264269
rect -50 -264343 50 -264327
rect -50 -264377 -34 -264343
rect 34 -264377 50 -264343
rect -50 -264415 50 -264377
rect -50 -265453 50 -265415
rect -50 -265487 -34 -265453
rect 34 -265487 50 -265453
rect -50 -265503 50 -265487
rect -50 -265561 50 -265545
rect -50 -265595 -34 -265561
rect 34 -265595 50 -265561
rect -50 -265633 50 -265595
rect -50 -266671 50 -266633
rect -50 -266705 -34 -266671
rect 34 -266705 50 -266671
rect -50 -266721 50 -266705
rect -50 -266779 50 -266763
rect -50 -266813 -34 -266779
rect 34 -266813 50 -266779
rect -50 -266851 50 -266813
rect -50 -267889 50 -267851
rect -50 -267923 -34 -267889
rect 34 -267923 50 -267889
rect -50 -267939 50 -267923
rect -50 -267997 50 -267981
rect -50 -268031 -34 -267997
rect 34 -268031 50 -267997
rect -50 -268069 50 -268031
rect -50 -269107 50 -269069
rect -50 -269141 -34 -269107
rect 34 -269141 50 -269107
rect -50 -269157 50 -269141
rect -50 -269215 50 -269199
rect -50 -269249 -34 -269215
rect 34 -269249 50 -269215
rect -50 -269287 50 -269249
rect -50 -270325 50 -270287
rect -50 -270359 -34 -270325
rect 34 -270359 50 -270325
rect -50 -270375 50 -270359
rect -50 -270433 50 -270417
rect -50 -270467 -34 -270433
rect 34 -270467 50 -270433
rect -50 -270505 50 -270467
rect -50 -271543 50 -271505
rect -50 -271577 -34 -271543
rect 34 -271577 50 -271543
rect -50 -271593 50 -271577
rect -50 -271651 50 -271635
rect -50 -271685 -34 -271651
rect 34 -271685 50 -271651
rect -50 -271723 50 -271685
rect -50 -272761 50 -272723
rect -50 -272795 -34 -272761
rect 34 -272795 50 -272761
rect -50 -272811 50 -272795
rect -50 -272869 50 -272853
rect -50 -272903 -34 -272869
rect 34 -272903 50 -272869
rect -50 -272941 50 -272903
rect -50 -273979 50 -273941
rect -50 -274013 -34 -273979
rect 34 -274013 50 -273979
rect -50 -274029 50 -274013
rect -50 -274087 50 -274071
rect -50 -274121 -34 -274087
rect 34 -274121 50 -274087
rect -50 -274159 50 -274121
rect -50 -275197 50 -275159
rect -50 -275231 -34 -275197
rect 34 -275231 50 -275197
rect -50 -275247 50 -275231
rect -50 -275305 50 -275289
rect -50 -275339 -34 -275305
rect 34 -275339 50 -275305
rect -50 -275377 50 -275339
rect -50 -276415 50 -276377
rect -50 -276449 -34 -276415
rect 34 -276449 50 -276415
rect -50 -276465 50 -276449
rect -50 -276523 50 -276507
rect -50 -276557 -34 -276523
rect 34 -276557 50 -276523
rect -50 -276595 50 -276557
rect -50 -277633 50 -277595
rect -50 -277667 -34 -277633
rect 34 -277667 50 -277633
rect -50 -277683 50 -277667
rect -50 -277741 50 -277725
rect -50 -277775 -34 -277741
rect 34 -277775 50 -277741
rect -50 -277813 50 -277775
rect -50 -278851 50 -278813
rect -50 -278885 -34 -278851
rect 34 -278885 50 -278851
rect -50 -278901 50 -278885
rect -50 -278959 50 -278943
rect -50 -278993 -34 -278959
rect 34 -278993 50 -278959
rect -50 -279031 50 -278993
rect -50 -280069 50 -280031
rect -50 -280103 -34 -280069
rect 34 -280103 50 -280069
rect -50 -280119 50 -280103
rect -50 -280177 50 -280161
rect -50 -280211 -34 -280177
rect 34 -280211 50 -280177
rect -50 -280249 50 -280211
rect -50 -281287 50 -281249
rect -50 -281321 -34 -281287
rect 34 -281321 50 -281287
rect -50 -281337 50 -281321
rect -50 -281395 50 -281379
rect -50 -281429 -34 -281395
rect 34 -281429 50 -281395
rect -50 -281467 50 -281429
rect -50 -282505 50 -282467
rect -50 -282539 -34 -282505
rect 34 -282539 50 -282505
rect -50 -282555 50 -282539
rect -50 -282613 50 -282597
rect -50 -282647 -34 -282613
rect 34 -282647 50 -282613
rect -50 -282685 50 -282647
rect -50 -283723 50 -283685
rect -50 -283757 -34 -283723
rect 34 -283757 50 -283723
rect -50 -283773 50 -283757
rect -50 -283831 50 -283815
rect -50 -283865 -34 -283831
rect 34 -283865 50 -283831
rect -50 -283903 50 -283865
rect -50 -284941 50 -284903
rect -50 -284975 -34 -284941
rect 34 -284975 50 -284941
rect -50 -284991 50 -284975
rect -50 -285049 50 -285033
rect -50 -285083 -34 -285049
rect 34 -285083 50 -285049
rect -50 -285121 50 -285083
rect -50 -286159 50 -286121
rect -50 -286193 -34 -286159
rect 34 -286193 50 -286159
rect -50 -286209 50 -286193
rect -50 -286267 50 -286251
rect -50 -286301 -34 -286267
rect 34 -286301 50 -286267
rect -50 -286339 50 -286301
rect -50 -287377 50 -287339
rect -50 -287411 -34 -287377
rect 34 -287411 50 -287377
rect -50 -287427 50 -287411
rect -50 -287485 50 -287469
rect -50 -287519 -34 -287485
rect 34 -287519 50 -287485
rect -50 -287557 50 -287519
rect -50 -288595 50 -288557
rect -50 -288629 -34 -288595
rect 34 -288629 50 -288595
rect -50 -288645 50 -288629
rect -50 -288703 50 -288687
rect -50 -288737 -34 -288703
rect 34 -288737 50 -288703
rect -50 -288775 50 -288737
rect -50 -289813 50 -289775
rect -50 -289847 -34 -289813
rect 34 -289847 50 -289813
rect -50 -289863 50 -289847
rect -50 -289921 50 -289905
rect -50 -289955 -34 -289921
rect 34 -289955 50 -289921
rect -50 -289993 50 -289955
rect -50 -291031 50 -290993
rect -50 -291065 -34 -291031
rect 34 -291065 50 -291031
rect -50 -291081 50 -291065
rect -50 -291139 50 -291123
rect -50 -291173 -34 -291139
rect 34 -291173 50 -291139
rect -50 -291211 50 -291173
rect -50 -292249 50 -292211
rect -50 -292283 -34 -292249
rect 34 -292283 50 -292249
rect -50 -292299 50 -292283
rect -50 -292357 50 -292341
rect -50 -292391 -34 -292357
rect 34 -292391 50 -292357
rect -50 -292429 50 -292391
rect -50 -293467 50 -293429
rect -50 -293501 -34 -293467
rect 34 -293501 50 -293467
rect -50 -293517 50 -293501
rect -50 -293575 50 -293559
rect -50 -293609 -34 -293575
rect 34 -293609 50 -293575
rect -50 -293647 50 -293609
rect -50 -294685 50 -294647
rect -50 -294719 -34 -294685
rect 34 -294719 50 -294685
rect -50 -294735 50 -294719
rect -50 -294793 50 -294777
rect -50 -294827 -34 -294793
rect 34 -294827 50 -294793
rect -50 -294865 50 -294827
rect -50 -295903 50 -295865
rect -50 -295937 -34 -295903
rect 34 -295937 50 -295903
rect -50 -295953 50 -295937
rect -50 -296011 50 -295995
rect -50 -296045 -34 -296011
rect 34 -296045 50 -296011
rect -50 -296083 50 -296045
rect -50 -297121 50 -297083
rect -50 -297155 -34 -297121
rect 34 -297155 50 -297121
rect -50 -297171 50 -297155
rect -50 -297229 50 -297213
rect -50 -297263 -34 -297229
rect 34 -297263 50 -297229
rect -50 -297301 50 -297263
rect -50 -298339 50 -298301
rect -50 -298373 -34 -298339
rect 34 -298373 50 -298339
rect -50 -298389 50 -298373
rect -50 -298447 50 -298431
rect -50 -298481 -34 -298447
rect 34 -298481 50 -298447
rect -50 -298519 50 -298481
rect -50 -299557 50 -299519
rect -50 -299591 -34 -299557
rect 34 -299591 50 -299557
rect -50 -299607 50 -299591
rect -50 -299665 50 -299649
rect -50 -299699 -34 -299665
rect 34 -299699 50 -299665
rect -50 -299737 50 -299699
rect -50 -300775 50 -300737
rect -50 -300809 -34 -300775
rect 34 -300809 50 -300775
rect -50 -300825 50 -300809
rect -50 -300883 50 -300867
rect -50 -300917 -34 -300883
rect 34 -300917 50 -300883
rect -50 -300955 50 -300917
rect -50 -301993 50 -301955
rect -50 -302027 -34 -301993
rect 34 -302027 50 -301993
rect -50 -302043 50 -302027
rect -50 -302101 50 -302085
rect -50 -302135 -34 -302101
rect 34 -302135 50 -302101
rect -50 -302173 50 -302135
rect -50 -303211 50 -303173
rect -50 -303245 -34 -303211
rect 34 -303245 50 -303211
rect -50 -303261 50 -303245
rect -50 -303319 50 -303303
rect -50 -303353 -34 -303319
rect 34 -303353 50 -303319
rect -50 -303391 50 -303353
rect -50 -304429 50 -304391
rect -50 -304463 -34 -304429
rect 34 -304463 50 -304429
rect -50 -304479 50 -304463
rect -50 -304537 50 -304521
rect -50 -304571 -34 -304537
rect 34 -304571 50 -304537
rect -50 -304609 50 -304571
rect -50 -305647 50 -305609
rect -50 -305681 -34 -305647
rect 34 -305681 50 -305647
rect -50 -305697 50 -305681
rect -50 -305755 50 -305739
rect -50 -305789 -34 -305755
rect 34 -305789 50 -305755
rect -50 -305827 50 -305789
rect -50 -306865 50 -306827
rect -50 -306899 -34 -306865
rect 34 -306899 50 -306865
rect -50 -306915 50 -306899
rect -50 -306973 50 -306957
rect -50 -307007 -34 -306973
rect 34 -307007 50 -306973
rect -50 -307045 50 -307007
rect -50 -308083 50 -308045
rect -50 -308117 -34 -308083
rect 34 -308117 50 -308083
rect -50 -308133 50 -308117
rect -50 -308191 50 -308175
rect -50 -308225 -34 -308191
rect 34 -308225 50 -308191
rect -50 -308263 50 -308225
rect -50 -309301 50 -309263
rect -50 -309335 -34 -309301
rect 34 -309335 50 -309301
rect -50 -309351 50 -309335
rect -50 -309409 50 -309393
rect -50 -309443 -34 -309409
rect 34 -309443 50 -309409
rect -50 -309481 50 -309443
rect -50 -310519 50 -310481
rect -50 -310553 -34 -310519
rect 34 -310553 50 -310519
rect -50 -310569 50 -310553
rect -50 -310627 50 -310611
rect -50 -310661 -34 -310627
rect 34 -310661 50 -310627
rect -50 -310699 50 -310661
rect -50 -311737 50 -311699
rect -50 -311771 -34 -311737
rect 34 -311771 50 -311737
rect -50 -311787 50 -311771
rect -50 -311845 50 -311829
rect -50 -311879 -34 -311845
rect 34 -311879 50 -311845
rect -50 -311917 50 -311879
rect -50 -312955 50 -312917
rect -50 -312989 -34 -312955
rect 34 -312989 50 -312955
rect -50 -313005 50 -312989
rect -50 -313063 50 -313047
rect -50 -313097 -34 -313063
rect 34 -313097 50 -313063
rect -50 -313135 50 -313097
rect -50 -314173 50 -314135
rect -50 -314207 -34 -314173
rect 34 -314207 50 -314173
rect -50 -314223 50 -314207
rect -50 -314281 50 -314265
rect -50 -314315 -34 -314281
rect 34 -314315 50 -314281
rect -50 -314353 50 -314315
rect -50 -315391 50 -315353
rect -50 -315425 -34 -315391
rect 34 -315425 50 -315391
rect -50 -315441 50 -315425
rect -50 -315499 50 -315483
rect -50 -315533 -34 -315499
rect 34 -315533 50 -315499
rect -50 -315571 50 -315533
rect -50 -316609 50 -316571
rect -50 -316643 -34 -316609
rect 34 -316643 50 -316609
rect -50 -316659 50 -316643
rect -50 -316717 50 -316701
rect -50 -316751 -34 -316717
rect 34 -316751 50 -316717
rect -50 -316789 50 -316751
rect -50 -317827 50 -317789
rect -50 -317861 -34 -317827
rect 34 -317861 50 -317827
rect -50 -317877 50 -317861
rect -50 -317935 50 -317919
rect -50 -317969 -34 -317935
rect 34 -317969 50 -317935
rect -50 -318007 50 -317969
rect -50 -319045 50 -319007
rect -50 -319079 -34 -319045
rect 34 -319079 50 -319045
rect -50 -319095 50 -319079
rect -50 -319153 50 -319137
rect -50 -319187 -34 -319153
rect 34 -319187 50 -319153
rect -50 -319225 50 -319187
rect -50 -320263 50 -320225
rect -50 -320297 -34 -320263
rect 34 -320297 50 -320263
rect -50 -320313 50 -320297
rect -50 -320371 50 -320355
rect -50 -320405 -34 -320371
rect 34 -320405 50 -320371
rect -50 -320443 50 -320405
rect -50 -321481 50 -321443
rect -50 -321515 -34 -321481
rect 34 -321515 50 -321481
rect -50 -321531 50 -321515
rect -50 -321589 50 -321573
rect -50 -321623 -34 -321589
rect 34 -321623 50 -321589
rect -50 -321661 50 -321623
rect -50 -322699 50 -322661
rect -50 -322733 -34 -322699
rect 34 -322733 50 -322699
rect -50 -322749 50 -322733
rect -50 -322807 50 -322791
rect -50 -322841 -34 -322807
rect 34 -322841 50 -322807
rect -50 -322879 50 -322841
rect -50 -323917 50 -323879
rect -50 -323951 -34 -323917
rect 34 -323951 50 -323917
rect -50 -323967 50 -323951
rect -50 -324025 50 -324009
rect -50 -324059 -34 -324025
rect 34 -324059 50 -324025
rect -50 -324097 50 -324059
rect -50 -325135 50 -325097
rect -50 -325169 -34 -325135
rect 34 -325169 50 -325135
rect -50 -325185 50 -325169
rect -50 -325243 50 -325227
rect -50 -325277 -34 -325243
rect 34 -325277 50 -325243
rect -50 -325315 50 -325277
rect -50 -326353 50 -326315
rect -50 -326387 -34 -326353
rect 34 -326387 50 -326353
rect -50 -326403 50 -326387
rect -50 -326461 50 -326445
rect -50 -326495 -34 -326461
rect 34 -326495 50 -326461
rect -50 -326533 50 -326495
rect -50 -327571 50 -327533
rect -50 -327605 -34 -327571
rect 34 -327605 50 -327571
rect -50 -327621 50 -327605
rect -50 -327679 50 -327663
rect -50 -327713 -34 -327679
rect 34 -327713 50 -327679
rect -50 -327751 50 -327713
rect -50 -328789 50 -328751
rect -50 -328823 -34 -328789
rect 34 -328823 50 -328789
rect -50 -328839 50 -328823
rect -50 -328897 50 -328881
rect -50 -328931 -34 -328897
rect 34 -328931 50 -328897
rect -50 -328969 50 -328931
rect -50 -330007 50 -329969
rect -50 -330041 -34 -330007
rect 34 -330041 50 -330007
rect -50 -330057 50 -330041
rect -50 -330115 50 -330099
rect -50 -330149 -34 -330115
rect 34 -330149 50 -330115
rect -50 -330187 50 -330149
rect -50 -331225 50 -331187
rect -50 -331259 -34 -331225
rect 34 -331259 50 -331225
rect -50 -331275 50 -331259
rect -50 -331333 50 -331317
rect -50 -331367 -34 -331333
rect 34 -331367 50 -331333
rect -50 -331405 50 -331367
rect -50 -332443 50 -332405
rect -50 -332477 -34 -332443
rect 34 -332477 50 -332443
rect -50 -332493 50 -332477
rect -50 -332551 50 -332535
rect -50 -332585 -34 -332551
rect 34 -332585 50 -332551
rect -50 -332623 50 -332585
rect -50 -333661 50 -333623
rect -50 -333695 -34 -333661
rect 34 -333695 50 -333661
rect -50 -333711 50 -333695
rect -50 -333769 50 -333753
rect -50 -333803 -34 -333769
rect 34 -333803 50 -333769
rect -50 -333841 50 -333803
rect -50 -334879 50 -334841
rect -50 -334913 -34 -334879
rect 34 -334913 50 -334879
rect -50 -334929 50 -334913
rect -50 -334987 50 -334971
rect -50 -335021 -34 -334987
rect 34 -335021 50 -334987
rect -50 -335059 50 -335021
rect -50 -336097 50 -336059
rect -50 -336131 -34 -336097
rect 34 -336131 50 -336097
rect -50 -336147 50 -336131
rect -50 -336205 50 -336189
rect -50 -336239 -34 -336205
rect 34 -336239 50 -336205
rect -50 -336277 50 -336239
rect -50 -337315 50 -337277
rect -50 -337349 -34 -337315
rect 34 -337349 50 -337315
rect -50 -337365 50 -337349
rect -50 -337423 50 -337407
rect -50 -337457 -34 -337423
rect 34 -337457 50 -337423
rect -50 -337495 50 -337457
rect -50 -338533 50 -338495
rect -50 -338567 -34 -338533
rect 34 -338567 50 -338533
rect -50 -338583 50 -338567
rect -50 -338641 50 -338625
rect -50 -338675 -34 -338641
rect 34 -338675 50 -338641
rect -50 -338713 50 -338675
rect -50 -339751 50 -339713
rect -50 -339785 -34 -339751
rect 34 -339785 50 -339751
rect -50 -339801 50 -339785
rect -50 -339859 50 -339843
rect -50 -339893 -34 -339859
rect 34 -339893 50 -339859
rect -50 -339931 50 -339893
rect -50 -340969 50 -340931
rect -50 -341003 -34 -340969
rect 34 -341003 50 -340969
rect -50 -341019 50 -341003
rect -50 -341077 50 -341061
rect -50 -341111 -34 -341077
rect 34 -341111 50 -341077
rect -50 -341149 50 -341111
rect -50 -342187 50 -342149
rect -50 -342221 -34 -342187
rect 34 -342221 50 -342187
rect -50 -342237 50 -342221
rect -50 -342295 50 -342279
rect -50 -342329 -34 -342295
rect 34 -342329 50 -342295
rect -50 -342367 50 -342329
rect -50 -343405 50 -343367
rect -50 -343439 -34 -343405
rect 34 -343439 50 -343405
rect -50 -343455 50 -343439
rect -50 -343513 50 -343497
rect -50 -343547 -34 -343513
rect 34 -343547 50 -343513
rect -50 -343585 50 -343547
rect -50 -344623 50 -344585
rect -50 -344657 -34 -344623
rect 34 -344657 50 -344623
rect -50 -344673 50 -344657
rect -50 -344731 50 -344715
rect -50 -344765 -34 -344731
rect 34 -344765 50 -344731
rect -50 -344803 50 -344765
rect -50 -345841 50 -345803
rect -50 -345875 -34 -345841
rect 34 -345875 50 -345841
rect -50 -345891 50 -345875
rect -50 -345949 50 -345933
rect -50 -345983 -34 -345949
rect 34 -345983 50 -345949
rect -50 -346021 50 -345983
rect -50 -347059 50 -347021
rect -50 -347093 -34 -347059
rect 34 -347093 50 -347059
rect -50 -347109 50 -347093
rect -50 -347167 50 -347151
rect -50 -347201 -34 -347167
rect 34 -347201 50 -347167
rect -50 -347239 50 -347201
rect -50 -348277 50 -348239
rect -50 -348311 -34 -348277
rect 34 -348311 50 -348277
rect -50 -348327 50 -348311
rect -50 -348385 50 -348369
rect -50 -348419 -34 -348385
rect 34 -348419 50 -348385
rect -50 -348457 50 -348419
rect -50 -349495 50 -349457
rect -50 -349529 -34 -349495
rect 34 -349529 50 -349495
rect -50 -349545 50 -349529
rect -50 -349603 50 -349587
rect -50 -349637 -34 -349603
rect 34 -349637 50 -349603
rect -50 -349675 50 -349637
rect -50 -350713 50 -350675
rect -50 -350747 -34 -350713
rect 34 -350747 50 -350713
rect -50 -350763 50 -350747
rect -50 -350821 50 -350805
rect -50 -350855 -34 -350821
rect 34 -350855 50 -350821
rect -50 -350893 50 -350855
rect -50 -351931 50 -351893
rect -50 -351965 -34 -351931
rect 34 -351965 50 -351931
rect -50 -351981 50 -351965
rect -50 -352039 50 -352023
rect -50 -352073 -34 -352039
rect 34 -352073 50 -352039
rect -50 -352111 50 -352073
rect -50 -353149 50 -353111
rect -50 -353183 -34 -353149
rect 34 -353183 50 -353149
rect -50 -353199 50 -353183
rect -50 -353257 50 -353241
rect -50 -353291 -34 -353257
rect 34 -353291 50 -353257
rect -50 -353329 50 -353291
rect -50 -354367 50 -354329
rect -50 -354401 -34 -354367
rect 34 -354401 50 -354367
rect -50 -354417 50 -354401
rect -50 -354475 50 -354459
rect -50 -354509 -34 -354475
rect 34 -354509 50 -354475
rect -50 -354547 50 -354509
rect -50 -355585 50 -355547
rect -50 -355619 -34 -355585
rect 34 -355619 50 -355585
rect -50 -355635 50 -355619
rect -50 -355693 50 -355677
rect -50 -355727 -34 -355693
rect 34 -355727 50 -355693
rect -50 -355765 50 -355727
rect -50 -356803 50 -356765
rect -50 -356837 -34 -356803
rect 34 -356837 50 -356803
rect -50 -356853 50 -356837
rect -50 -356911 50 -356895
rect -50 -356945 -34 -356911
rect 34 -356945 50 -356911
rect -50 -356983 50 -356945
rect -50 -358021 50 -357983
rect -50 -358055 -34 -358021
rect 34 -358055 50 -358021
rect -50 -358071 50 -358055
rect -50 -358129 50 -358113
rect -50 -358163 -34 -358129
rect 34 -358163 50 -358129
rect -50 -358201 50 -358163
rect -50 -359239 50 -359201
rect -50 -359273 -34 -359239
rect 34 -359273 50 -359239
rect -50 -359289 50 -359273
rect -50 -359347 50 -359331
rect -50 -359381 -34 -359347
rect 34 -359381 50 -359347
rect -50 -359419 50 -359381
rect -50 -360457 50 -360419
rect -50 -360491 -34 -360457
rect 34 -360491 50 -360457
rect -50 -360507 50 -360491
rect -50 -360565 50 -360549
rect -50 -360599 -34 -360565
rect 34 -360599 50 -360565
rect -50 -360637 50 -360599
rect -50 -361675 50 -361637
rect -50 -361709 -34 -361675
rect 34 -361709 50 -361675
rect -50 -361725 50 -361709
rect -50 -361783 50 -361767
rect -50 -361817 -34 -361783
rect 34 -361817 50 -361783
rect -50 -361855 50 -361817
rect -50 -362893 50 -362855
rect -50 -362927 -34 -362893
rect 34 -362927 50 -362893
rect -50 -362943 50 -362927
rect -50 -363001 50 -362985
rect -50 -363035 -34 -363001
rect 34 -363035 50 -363001
rect -50 -363073 50 -363035
rect -50 -364111 50 -364073
rect -50 -364145 -34 -364111
rect 34 -364145 50 -364111
rect -50 -364161 50 -364145
rect -50 -364219 50 -364203
rect -50 -364253 -34 -364219
rect 34 -364253 50 -364219
rect -50 -364291 50 -364253
rect -50 -365329 50 -365291
rect -50 -365363 -34 -365329
rect 34 -365363 50 -365329
rect -50 -365379 50 -365363
rect -50 -365437 50 -365421
rect -50 -365471 -34 -365437
rect 34 -365471 50 -365437
rect -50 -365509 50 -365471
rect -50 -366547 50 -366509
rect -50 -366581 -34 -366547
rect 34 -366581 50 -366547
rect -50 -366597 50 -366581
rect -50 -366655 50 -366639
rect -50 -366689 -34 -366655
rect 34 -366689 50 -366655
rect -50 -366727 50 -366689
rect -50 -367765 50 -367727
rect -50 -367799 -34 -367765
rect 34 -367799 50 -367765
rect -50 -367815 50 -367799
rect -50 -367873 50 -367857
rect -50 -367907 -34 -367873
rect 34 -367907 50 -367873
rect -50 -367945 50 -367907
rect -50 -368983 50 -368945
rect -50 -369017 -34 -368983
rect 34 -369017 50 -368983
rect -50 -369033 50 -369017
rect -50 -369091 50 -369075
rect -50 -369125 -34 -369091
rect 34 -369125 50 -369091
rect -50 -369163 50 -369125
rect -50 -370201 50 -370163
rect -50 -370235 -34 -370201
rect 34 -370235 50 -370201
rect -50 -370251 50 -370235
rect -50 -370309 50 -370293
rect -50 -370343 -34 -370309
rect 34 -370343 50 -370309
rect -50 -370381 50 -370343
rect -50 -371419 50 -371381
rect -50 -371453 -34 -371419
rect 34 -371453 50 -371419
rect -50 -371469 50 -371453
rect -50 -371527 50 -371511
rect -50 -371561 -34 -371527
rect 34 -371561 50 -371527
rect -50 -371599 50 -371561
rect -50 -372637 50 -372599
rect -50 -372671 -34 -372637
rect 34 -372671 50 -372637
rect -50 -372687 50 -372671
rect -50 -372745 50 -372729
rect -50 -372779 -34 -372745
rect 34 -372779 50 -372745
rect -50 -372817 50 -372779
rect -50 -373855 50 -373817
rect -50 -373889 -34 -373855
rect 34 -373889 50 -373855
rect -50 -373905 50 -373889
rect -50 -373963 50 -373947
rect -50 -373997 -34 -373963
rect 34 -373997 50 -373963
rect -50 -374035 50 -373997
rect -50 -375073 50 -375035
rect -50 -375107 -34 -375073
rect 34 -375107 50 -375073
rect -50 -375123 50 -375107
rect -50 -375181 50 -375165
rect -50 -375215 -34 -375181
rect 34 -375215 50 -375181
rect -50 -375253 50 -375215
rect -50 -376291 50 -376253
rect -50 -376325 -34 -376291
rect 34 -376325 50 -376291
rect -50 -376341 50 -376325
rect -50 -376399 50 -376383
rect -50 -376433 -34 -376399
rect 34 -376433 50 -376399
rect -50 -376471 50 -376433
rect -50 -377509 50 -377471
rect -50 -377543 -34 -377509
rect 34 -377543 50 -377509
rect -50 -377559 50 -377543
rect -50 -377617 50 -377601
rect -50 -377651 -34 -377617
rect 34 -377651 50 -377617
rect -50 -377689 50 -377651
rect -50 -378727 50 -378689
rect -50 -378761 -34 -378727
rect 34 -378761 50 -378727
rect -50 -378777 50 -378761
rect -50 -378835 50 -378819
rect -50 -378869 -34 -378835
rect 34 -378869 50 -378835
rect -50 -378907 50 -378869
rect -50 -379945 50 -379907
rect -50 -379979 -34 -379945
rect 34 -379979 50 -379945
rect -50 -379995 50 -379979
rect -50 -380053 50 -380037
rect -50 -380087 -34 -380053
rect 34 -380087 50 -380053
rect -50 -380125 50 -380087
rect -50 -381163 50 -381125
rect -50 -381197 -34 -381163
rect 34 -381197 50 -381163
rect -50 -381213 50 -381197
rect -50 -381271 50 -381255
rect -50 -381305 -34 -381271
rect 34 -381305 50 -381271
rect -50 -381343 50 -381305
rect -50 -382381 50 -382343
rect -50 -382415 -34 -382381
rect 34 -382415 50 -382381
rect -50 -382431 50 -382415
rect -50 -382489 50 -382473
rect -50 -382523 -34 -382489
rect 34 -382523 50 -382489
rect -50 -382561 50 -382523
rect -50 -383599 50 -383561
rect -50 -383633 -34 -383599
rect 34 -383633 50 -383599
rect -50 -383649 50 -383633
rect -50 -383707 50 -383691
rect -50 -383741 -34 -383707
rect 34 -383741 50 -383707
rect -50 -383779 50 -383741
rect -50 -384817 50 -384779
rect -50 -384851 -34 -384817
rect 34 -384851 50 -384817
rect -50 -384867 50 -384851
rect -50 -384925 50 -384909
rect -50 -384959 -34 -384925
rect 34 -384959 50 -384925
rect -50 -384997 50 -384959
rect -50 -386035 50 -385997
rect -50 -386069 -34 -386035
rect 34 -386069 50 -386035
rect -50 -386085 50 -386069
rect -50 -386143 50 -386127
rect -50 -386177 -34 -386143
rect 34 -386177 50 -386143
rect -50 -386215 50 -386177
rect -50 -387253 50 -387215
rect -50 -387287 -34 -387253
rect 34 -387287 50 -387253
rect -50 -387303 50 -387287
rect -50 -387361 50 -387345
rect -50 -387395 -34 -387361
rect 34 -387395 50 -387361
rect -50 -387433 50 -387395
rect -50 -388471 50 -388433
rect -50 -388505 -34 -388471
rect 34 -388505 50 -388471
rect -50 -388521 50 -388505
rect -50 -388579 50 -388563
rect -50 -388613 -34 -388579
rect 34 -388613 50 -388579
rect -50 -388651 50 -388613
rect -50 -389689 50 -389651
rect -50 -389723 -34 -389689
rect 34 -389723 50 -389689
rect -50 -389739 50 -389723
rect -50 -389797 50 -389781
rect -50 -389831 -34 -389797
rect 34 -389831 50 -389797
rect -50 -389869 50 -389831
rect -50 -390907 50 -390869
rect -50 -390941 -34 -390907
rect 34 -390941 50 -390907
rect -50 -390957 50 -390941
rect -50 -391015 50 -390999
rect -50 -391049 -34 -391015
rect 34 -391049 50 -391015
rect -50 -391087 50 -391049
rect -50 -392125 50 -392087
rect -50 -392159 -34 -392125
rect 34 -392159 50 -392125
rect -50 -392175 50 -392159
rect -50 -392233 50 -392217
rect -50 -392267 -34 -392233
rect 34 -392267 50 -392233
rect -50 -392305 50 -392267
rect -50 -393343 50 -393305
rect -50 -393377 -34 -393343
rect 34 -393377 50 -393343
rect -50 -393393 50 -393377
rect -50 -393451 50 -393435
rect -50 -393485 -34 -393451
rect 34 -393485 50 -393451
rect -50 -393523 50 -393485
rect -50 -394561 50 -394523
rect -50 -394595 -34 -394561
rect 34 -394595 50 -394561
rect -50 -394611 50 -394595
rect -50 -394669 50 -394653
rect -50 -394703 -34 -394669
rect 34 -394703 50 -394669
rect -50 -394741 50 -394703
rect -50 -395779 50 -395741
rect -50 -395813 -34 -395779
rect 34 -395813 50 -395779
rect -50 -395829 50 -395813
rect -50 -395887 50 -395871
rect -50 -395921 -34 -395887
rect 34 -395921 50 -395887
rect -50 -395959 50 -395921
rect -50 -396997 50 -396959
rect -50 -397031 -34 -396997
rect 34 -397031 50 -396997
rect -50 -397047 50 -397031
rect -50 -397105 50 -397089
rect -50 -397139 -34 -397105
rect 34 -397139 50 -397105
rect -50 -397177 50 -397139
rect -50 -398215 50 -398177
rect -50 -398249 -34 -398215
rect 34 -398249 50 -398215
rect -50 -398265 50 -398249
rect -50 -398323 50 -398307
rect -50 -398357 -34 -398323
rect 34 -398357 50 -398323
rect -50 -398395 50 -398357
rect -50 -399433 50 -399395
rect -50 -399467 -34 -399433
rect 34 -399467 50 -399433
rect -50 -399483 50 -399467
rect -50 -399541 50 -399525
rect -50 -399575 -34 -399541
rect 34 -399575 50 -399541
rect -50 -399613 50 -399575
rect -50 -400651 50 -400613
rect -50 -400685 -34 -400651
rect 34 -400685 50 -400651
rect -50 -400701 50 -400685
rect -50 -400759 50 -400743
rect -50 -400793 -34 -400759
rect 34 -400793 50 -400759
rect -50 -400831 50 -400793
rect -50 -401869 50 -401831
rect -50 -401903 -34 -401869
rect 34 -401903 50 -401869
rect -50 -401919 50 -401903
rect -50 -401977 50 -401961
rect -50 -402011 -34 -401977
rect 34 -402011 50 -401977
rect -50 -402049 50 -402011
rect -50 -403087 50 -403049
rect -50 -403121 -34 -403087
rect 34 -403121 50 -403087
rect -50 -403137 50 -403121
rect -50 -403195 50 -403179
rect -50 -403229 -34 -403195
rect 34 -403229 50 -403195
rect -50 -403267 50 -403229
rect -50 -404305 50 -404267
rect -50 -404339 -34 -404305
rect 34 -404339 50 -404305
rect -50 -404355 50 -404339
rect -50 -404413 50 -404397
rect -50 -404447 -34 -404413
rect 34 -404447 50 -404413
rect -50 -404485 50 -404447
rect -50 -405523 50 -405485
rect -50 -405557 -34 -405523
rect 34 -405557 50 -405523
rect -50 -405573 50 -405557
rect -50 -405631 50 -405615
rect -50 -405665 -34 -405631
rect 34 -405665 50 -405631
rect -50 -405703 50 -405665
rect -50 -406741 50 -406703
rect -50 -406775 -34 -406741
rect 34 -406775 50 -406741
rect -50 -406791 50 -406775
rect -50 -406849 50 -406833
rect -50 -406883 -34 -406849
rect 34 -406883 50 -406849
rect -50 -406921 50 -406883
rect -50 -407959 50 -407921
rect -50 -407993 -34 -407959
rect 34 -407993 50 -407959
rect -50 -408009 50 -407993
rect -50 -408067 50 -408051
rect -50 -408101 -34 -408067
rect 34 -408101 50 -408067
rect -50 -408139 50 -408101
rect -50 -409177 50 -409139
rect -50 -409211 -34 -409177
rect 34 -409211 50 -409177
rect -50 -409227 50 -409211
rect -50 -409285 50 -409269
rect -50 -409319 -34 -409285
rect 34 -409319 50 -409285
rect -50 -409357 50 -409319
rect -50 -410395 50 -410357
rect -50 -410429 -34 -410395
rect 34 -410429 50 -410395
rect -50 -410445 50 -410429
rect -50 -410503 50 -410487
rect -50 -410537 -34 -410503
rect 34 -410537 50 -410503
rect -50 -410575 50 -410537
rect -50 -411613 50 -411575
rect -50 -411647 -34 -411613
rect 34 -411647 50 -411613
rect -50 -411663 50 -411647
rect -50 -411721 50 -411705
rect -50 -411755 -34 -411721
rect 34 -411755 50 -411721
rect -50 -411793 50 -411755
rect -50 -412831 50 -412793
rect -50 -412865 -34 -412831
rect 34 -412865 50 -412831
rect -50 -412881 50 -412865
rect -50 -412939 50 -412923
rect -50 -412973 -34 -412939
rect 34 -412973 50 -412939
rect -50 -413011 50 -412973
rect -50 -414049 50 -414011
rect -50 -414083 -34 -414049
rect 34 -414083 50 -414049
rect -50 -414099 50 -414083
rect -50 -414157 50 -414141
rect -50 -414191 -34 -414157
rect 34 -414191 50 -414157
rect -50 -414229 50 -414191
rect -50 -415267 50 -415229
rect -50 -415301 -34 -415267
rect 34 -415301 50 -415267
rect -50 -415317 50 -415301
rect -50 -415375 50 -415359
rect -50 -415409 -34 -415375
rect 34 -415409 50 -415375
rect -50 -415447 50 -415409
rect -50 -416485 50 -416447
rect -50 -416519 -34 -416485
rect 34 -416519 50 -416485
rect -50 -416535 50 -416519
rect -50 -416593 50 -416577
rect -50 -416627 -34 -416593
rect 34 -416627 50 -416593
rect -50 -416665 50 -416627
rect -50 -417703 50 -417665
rect -50 -417737 -34 -417703
rect 34 -417737 50 -417703
rect -50 -417753 50 -417737
rect -50 -417811 50 -417795
rect -50 -417845 -34 -417811
rect 34 -417845 50 -417811
rect -50 -417883 50 -417845
rect -50 -418921 50 -418883
rect -50 -418955 -34 -418921
rect 34 -418955 50 -418921
rect -50 -418971 50 -418955
rect -50 -419029 50 -419013
rect -50 -419063 -34 -419029
rect 34 -419063 50 -419029
rect -50 -419101 50 -419063
rect -50 -420139 50 -420101
rect -50 -420173 -34 -420139
rect 34 -420173 50 -420139
rect -50 -420189 50 -420173
rect -50 -420247 50 -420231
rect -50 -420281 -34 -420247
rect 34 -420281 50 -420247
rect -50 -420319 50 -420281
rect -50 -421357 50 -421319
rect -50 -421391 -34 -421357
rect 34 -421391 50 -421357
rect -50 -421407 50 -421391
rect -50 -421465 50 -421449
rect -50 -421499 -34 -421465
rect 34 -421499 50 -421465
rect -50 -421537 50 -421499
rect -50 -422575 50 -422537
rect -50 -422609 -34 -422575
rect 34 -422609 50 -422575
rect -50 -422625 50 -422609
rect -50 -422683 50 -422667
rect -50 -422717 -34 -422683
rect 34 -422717 50 -422683
rect -50 -422755 50 -422717
rect -50 -423793 50 -423755
rect -50 -423827 -34 -423793
rect 34 -423827 50 -423793
rect -50 -423843 50 -423827
rect -50 -423901 50 -423885
rect -50 -423935 -34 -423901
rect 34 -423935 50 -423901
rect -50 -423973 50 -423935
rect -50 -425011 50 -424973
rect -50 -425045 -34 -425011
rect 34 -425045 50 -425011
rect -50 -425061 50 -425045
rect -50 -425119 50 -425103
rect -50 -425153 -34 -425119
rect 34 -425153 50 -425119
rect -50 -425191 50 -425153
rect -50 -426229 50 -426191
rect -50 -426263 -34 -426229
rect 34 -426263 50 -426229
rect -50 -426279 50 -426263
rect -50 -426337 50 -426321
rect -50 -426371 -34 -426337
rect 34 -426371 50 -426337
rect -50 -426409 50 -426371
rect -50 -427447 50 -427409
rect -50 -427481 -34 -427447
rect 34 -427481 50 -427447
rect -50 -427497 50 -427481
rect -50 -427555 50 -427539
rect -50 -427589 -34 -427555
rect 34 -427589 50 -427555
rect -50 -427627 50 -427589
rect -50 -428665 50 -428627
rect -50 -428699 -34 -428665
rect 34 -428699 50 -428665
rect -50 -428715 50 -428699
rect -50 -428773 50 -428757
rect -50 -428807 -34 -428773
rect 34 -428807 50 -428773
rect -50 -428845 50 -428807
rect -50 -429883 50 -429845
rect -50 -429917 -34 -429883
rect 34 -429917 50 -429883
rect -50 -429933 50 -429917
rect -50 -429991 50 -429975
rect -50 -430025 -34 -429991
rect 34 -430025 50 -429991
rect -50 -430063 50 -430025
rect -50 -431101 50 -431063
rect -50 -431135 -34 -431101
rect 34 -431135 50 -431101
rect -50 -431151 50 -431135
rect -50 -431209 50 -431193
rect -50 -431243 -34 -431209
rect 34 -431243 50 -431209
rect -50 -431281 50 -431243
rect -50 -432319 50 -432281
rect -50 -432353 -34 -432319
rect 34 -432353 50 -432319
rect -50 -432369 50 -432353
rect -50 -432427 50 -432411
rect -50 -432461 -34 -432427
rect 34 -432461 50 -432427
rect -50 -432499 50 -432461
rect -50 -433537 50 -433499
rect -50 -433571 -34 -433537
rect 34 -433571 50 -433537
rect -50 -433587 50 -433571
rect -50 -433645 50 -433629
rect -50 -433679 -34 -433645
rect 34 -433679 50 -433645
rect -50 -433717 50 -433679
rect -50 -434755 50 -434717
rect -50 -434789 -34 -434755
rect 34 -434789 50 -434755
rect -50 -434805 50 -434789
rect -50 -434863 50 -434847
rect -50 -434897 -34 -434863
rect 34 -434897 50 -434863
rect -50 -434935 50 -434897
rect -50 -435973 50 -435935
rect -50 -436007 -34 -435973
rect 34 -436007 50 -435973
rect -50 -436023 50 -436007
rect -50 -436081 50 -436065
rect -50 -436115 -34 -436081
rect 34 -436115 50 -436081
rect -50 -436153 50 -436115
rect -50 -437191 50 -437153
rect -50 -437225 -34 -437191
rect 34 -437225 50 -437191
rect -50 -437241 50 -437225
rect -50 -437299 50 -437283
rect -50 -437333 -34 -437299
rect 34 -437333 50 -437299
rect -50 -437371 50 -437333
rect -50 -438409 50 -438371
rect -50 -438443 -34 -438409
rect 34 -438443 50 -438409
rect -50 -438459 50 -438443
rect -50 -438517 50 -438501
rect -50 -438551 -34 -438517
rect 34 -438551 50 -438517
rect -50 -438589 50 -438551
rect -50 -439627 50 -439589
rect -50 -439661 -34 -439627
rect 34 -439661 50 -439627
rect -50 -439677 50 -439661
rect -50 -439735 50 -439719
rect -50 -439769 -34 -439735
rect 34 -439769 50 -439735
rect -50 -439807 50 -439769
rect -50 -440845 50 -440807
rect -50 -440879 -34 -440845
rect 34 -440879 50 -440845
rect -50 -440895 50 -440879
rect -50 -440953 50 -440937
rect -50 -440987 -34 -440953
rect 34 -440987 50 -440953
rect -50 -441025 50 -440987
rect -50 -442063 50 -442025
rect -50 -442097 -34 -442063
rect 34 -442097 50 -442063
rect -50 -442113 50 -442097
rect -50 -442171 50 -442155
rect -50 -442205 -34 -442171
rect 34 -442205 50 -442171
rect -50 -442243 50 -442205
rect -50 -443281 50 -443243
rect -50 -443315 -34 -443281
rect 34 -443315 50 -443281
rect -50 -443331 50 -443315
rect -50 -443389 50 -443373
rect -50 -443423 -34 -443389
rect 34 -443423 50 -443389
rect -50 -443461 50 -443423
rect -50 -444499 50 -444461
rect -50 -444533 -34 -444499
rect 34 -444533 50 -444499
rect -50 -444549 50 -444533
rect -50 -444607 50 -444591
rect -50 -444641 -34 -444607
rect 34 -444641 50 -444607
rect -50 -444679 50 -444641
rect -50 -445717 50 -445679
rect -50 -445751 -34 -445717
rect 34 -445751 50 -445717
rect -50 -445767 50 -445751
rect -50 -445825 50 -445809
rect -50 -445859 -34 -445825
rect 34 -445859 50 -445825
rect -50 -445897 50 -445859
rect -50 -446935 50 -446897
rect -50 -446969 -34 -446935
rect 34 -446969 50 -446935
rect -50 -446985 50 -446969
rect -50 -447043 50 -447027
rect -50 -447077 -34 -447043
rect 34 -447077 50 -447043
rect -50 -447115 50 -447077
rect -50 -448153 50 -448115
rect -50 -448187 -34 -448153
rect 34 -448187 50 -448153
rect -50 -448203 50 -448187
rect -50 -448261 50 -448245
rect -50 -448295 -34 -448261
rect 34 -448295 50 -448261
rect -50 -448333 50 -448295
rect -50 -449371 50 -449333
rect -50 -449405 -34 -449371
rect 34 -449405 50 -449371
rect -50 -449421 50 -449405
rect -50 -449479 50 -449463
rect -50 -449513 -34 -449479
rect 34 -449513 50 -449479
rect -50 -449551 50 -449513
rect -50 -450589 50 -450551
rect -50 -450623 -34 -450589
rect 34 -450623 50 -450589
rect -50 -450639 50 -450623
rect -50 -450697 50 -450681
rect -50 -450731 -34 -450697
rect 34 -450731 50 -450697
rect -50 -450769 50 -450731
rect -50 -451807 50 -451769
rect -50 -451841 -34 -451807
rect 34 -451841 50 -451807
rect -50 -451857 50 -451841
rect -50 -451915 50 -451899
rect -50 -451949 -34 -451915
rect 34 -451949 50 -451915
rect -50 -451987 50 -451949
rect -50 -453025 50 -452987
rect -50 -453059 -34 -453025
rect 34 -453059 50 -453025
rect -50 -453075 50 -453059
rect -50 -453133 50 -453117
rect -50 -453167 -34 -453133
rect 34 -453167 50 -453133
rect -50 -453205 50 -453167
rect -50 -454243 50 -454205
rect -50 -454277 -34 -454243
rect 34 -454277 50 -454243
rect -50 -454293 50 -454277
rect -50 -454351 50 -454335
rect -50 -454385 -34 -454351
rect 34 -454385 50 -454351
rect -50 -454423 50 -454385
rect -50 -455461 50 -455423
rect -50 -455495 -34 -455461
rect 34 -455495 50 -455461
rect -50 -455511 50 -455495
rect -50 -455569 50 -455553
rect -50 -455603 -34 -455569
rect 34 -455603 50 -455569
rect -50 -455641 50 -455603
rect -50 -456679 50 -456641
rect -50 -456713 -34 -456679
rect 34 -456713 50 -456679
rect -50 -456729 50 -456713
rect -50 -456787 50 -456771
rect -50 -456821 -34 -456787
rect 34 -456821 50 -456787
rect -50 -456859 50 -456821
rect -50 -457897 50 -457859
rect -50 -457931 -34 -457897
rect 34 -457931 50 -457897
rect -50 -457947 50 -457931
rect -50 -458005 50 -457989
rect -50 -458039 -34 -458005
rect 34 -458039 50 -458005
rect -50 -458077 50 -458039
rect -50 -459115 50 -459077
rect -50 -459149 -34 -459115
rect 34 -459149 50 -459115
rect -50 -459165 50 -459149
rect -50 -459223 50 -459207
rect -50 -459257 -34 -459223
rect 34 -459257 50 -459223
rect -50 -459295 50 -459257
rect -50 -460333 50 -460295
rect -50 -460367 -34 -460333
rect 34 -460367 50 -460333
rect -50 -460383 50 -460367
rect -50 -460441 50 -460425
rect -50 -460475 -34 -460441
rect 34 -460475 50 -460441
rect -50 -460513 50 -460475
rect -50 -461551 50 -461513
rect -50 -461585 -34 -461551
rect 34 -461585 50 -461551
rect -50 -461601 50 -461585
rect -50 -461659 50 -461643
rect -50 -461693 -34 -461659
rect 34 -461693 50 -461659
rect -50 -461731 50 -461693
rect -50 -462769 50 -462731
rect -50 -462803 -34 -462769
rect 34 -462803 50 -462769
rect -50 -462819 50 -462803
rect -50 -462877 50 -462861
rect -50 -462911 -34 -462877
rect 34 -462911 50 -462877
rect -50 -462949 50 -462911
rect -50 -463987 50 -463949
rect -50 -464021 -34 -463987
rect 34 -464021 50 -463987
rect -50 -464037 50 -464021
rect -50 -464095 50 -464079
rect -50 -464129 -34 -464095
rect 34 -464129 50 -464095
rect -50 -464167 50 -464129
rect -50 -465205 50 -465167
rect -50 -465239 -34 -465205
rect 34 -465239 50 -465205
rect -50 -465255 50 -465239
rect -50 -465313 50 -465297
rect -50 -465347 -34 -465313
rect 34 -465347 50 -465313
rect -50 -465385 50 -465347
rect -50 -466423 50 -466385
rect -50 -466457 -34 -466423
rect 34 -466457 50 -466423
rect -50 -466473 50 -466457
rect -50 -466531 50 -466515
rect -50 -466565 -34 -466531
rect 34 -466565 50 -466531
rect -50 -466603 50 -466565
rect -50 -467641 50 -467603
rect -50 -467675 -34 -467641
rect 34 -467675 50 -467641
rect -50 -467691 50 -467675
rect -50 -467749 50 -467733
rect -50 -467783 -34 -467749
rect 34 -467783 50 -467749
rect -50 -467821 50 -467783
rect -50 -468859 50 -468821
rect -50 -468893 -34 -468859
rect 34 -468893 50 -468859
rect -50 -468909 50 -468893
rect -50 -468967 50 -468951
rect -50 -469001 -34 -468967
rect 34 -469001 50 -468967
rect -50 -469039 50 -469001
rect -50 -470077 50 -470039
rect -50 -470111 -34 -470077
rect 34 -470111 50 -470077
rect -50 -470127 50 -470111
rect -50 -470185 50 -470169
rect -50 -470219 -34 -470185
rect 34 -470219 50 -470185
rect -50 -470257 50 -470219
rect -50 -471295 50 -471257
rect -50 -471329 -34 -471295
rect 34 -471329 50 -471295
rect -50 -471345 50 -471329
rect -50 -471403 50 -471387
rect -50 -471437 -34 -471403
rect 34 -471437 50 -471403
rect -50 -471475 50 -471437
rect -50 -472513 50 -472475
rect -50 -472547 -34 -472513
rect 34 -472547 50 -472513
rect -50 -472563 50 -472547
rect -50 -472621 50 -472605
rect -50 -472655 -34 -472621
rect 34 -472655 50 -472621
rect -50 -472693 50 -472655
rect -50 -473731 50 -473693
rect -50 -473765 -34 -473731
rect 34 -473765 50 -473731
rect -50 -473781 50 -473765
rect -50 -473839 50 -473823
rect -50 -473873 -34 -473839
rect 34 -473873 50 -473839
rect -50 -473911 50 -473873
rect -50 -474949 50 -474911
rect -50 -474983 -34 -474949
rect 34 -474983 50 -474949
rect -50 -474999 50 -474983
rect -50 -475057 50 -475041
rect -50 -475091 -34 -475057
rect 34 -475091 50 -475057
rect -50 -475129 50 -475091
rect -50 -476167 50 -476129
rect -50 -476201 -34 -476167
rect 34 -476201 50 -476167
rect -50 -476217 50 -476201
rect -50 -476275 50 -476259
rect -50 -476309 -34 -476275
rect 34 -476309 50 -476275
rect -50 -476347 50 -476309
rect -50 -477385 50 -477347
rect -50 -477419 -34 -477385
rect 34 -477419 50 -477385
rect -50 -477435 50 -477419
rect -50 -477493 50 -477477
rect -50 -477527 -34 -477493
rect 34 -477527 50 -477493
rect -50 -477565 50 -477527
rect -50 -478603 50 -478565
rect -50 -478637 -34 -478603
rect 34 -478637 50 -478603
rect -50 -478653 50 -478637
rect -50 -478711 50 -478695
rect -50 -478745 -34 -478711
rect 34 -478745 50 -478711
rect -50 -478783 50 -478745
rect -50 -479821 50 -479783
rect -50 -479855 -34 -479821
rect 34 -479855 50 -479821
rect -50 -479871 50 -479855
rect -50 -479929 50 -479913
rect -50 -479963 -34 -479929
rect 34 -479963 50 -479929
rect -50 -480001 50 -479963
rect -50 -481039 50 -481001
rect -50 -481073 -34 -481039
rect 34 -481073 50 -481039
rect -50 -481089 50 -481073
rect -50 -481147 50 -481131
rect -50 -481181 -34 -481147
rect 34 -481181 50 -481147
rect -50 -481219 50 -481181
rect -50 -482257 50 -482219
rect -50 -482291 -34 -482257
rect 34 -482291 50 -482257
rect -50 -482307 50 -482291
rect -50 -482365 50 -482349
rect -50 -482399 -34 -482365
rect 34 -482399 50 -482365
rect -50 -482437 50 -482399
rect -50 -483475 50 -483437
rect -50 -483509 -34 -483475
rect 34 -483509 50 -483475
rect -50 -483525 50 -483509
rect -50 -483583 50 -483567
rect -50 -483617 -34 -483583
rect 34 -483617 50 -483583
rect -50 -483655 50 -483617
rect -50 -484693 50 -484655
rect -50 -484727 -34 -484693
rect 34 -484727 50 -484693
rect -50 -484743 50 -484727
rect -50 -484801 50 -484785
rect -50 -484835 -34 -484801
rect 34 -484835 50 -484801
rect -50 -484873 50 -484835
rect -50 -485911 50 -485873
rect -50 -485945 -34 -485911
rect 34 -485945 50 -485911
rect -50 -485961 50 -485945
rect -50 -486019 50 -486003
rect -50 -486053 -34 -486019
rect 34 -486053 50 -486019
rect -50 -486091 50 -486053
rect -50 -487129 50 -487091
rect -50 -487163 -34 -487129
rect 34 -487163 50 -487129
rect -50 -487179 50 -487163
rect -50 -487237 50 -487221
rect -50 -487271 -34 -487237
rect 34 -487271 50 -487237
rect -50 -487309 50 -487271
rect -50 -488347 50 -488309
rect -50 -488381 -34 -488347
rect 34 -488381 50 -488347
rect -50 -488397 50 -488381
rect -50 -488455 50 -488439
rect -50 -488489 -34 -488455
rect 34 -488489 50 -488455
rect -50 -488527 50 -488489
rect -50 -489565 50 -489527
rect -50 -489599 -34 -489565
rect 34 -489599 50 -489565
rect -50 -489615 50 -489599
rect -50 -489673 50 -489657
rect -50 -489707 -34 -489673
rect 34 -489707 50 -489673
rect -50 -489745 50 -489707
rect -50 -490783 50 -490745
rect -50 -490817 -34 -490783
rect 34 -490817 50 -490783
rect -50 -490833 50 -490817
rect -50 -490891 50 -490875
rect -50 -490925 -34 -490891
rect 34 -490925 50 -490891
rect -50 -490963 50 -490925
rect -50 -492001 50 -491963
rect -50 -492035 -34 -492001
rect 34 -492035 50 -492001
rect -50 -492051 50 -492035
rect -50 -492109 50 -492093
rect -50 -492143 -34 -492109
rect 34 -492143 50 -492109
rect -50 -492181 50 -492143
rect -50 -493219 50 -493181
rect -50 -493253 -34 -493219
rect 34 -493253 50 -493219
rect -50 -493269 50 -493253
rect -50 -493327 50 -493311
rect -50 -493361 -34 -493327
rect 34 -493361 50 -493327
rect -50 -493399 50 -493361
rect -50 -494437 50 -494399
rect -50 -494471 -34 -494437
rect 34 -494471 50 -494437
rect -50 -494487 50 -494471
rect -50 -494545 50 -494529
rect -50 -494579 -34 -494545
rect 34 -494579 50 -494545
rect -50 -494617 50 -494579
rect -50 -495655 50 -495617
rect -50 -495689 -34 -495655
rect 34 -495689 50 -495655
rect -50 -495705 50 -495689
rect -50 -495763 50 -495747
rect -50 -495797 -34 -495763
rect 34 -495797 50 -495763
rect -50 -495835 50 -495797
rect -50 -496873 50 -496835
rect -50 -496907 -34 -496873
rect 34 -496907 50 -496873
rect -50 -496923 50 -496907
rect -50 -496981 50 -496965
rect -50 -497015 -34 -496981
rect 34 -497015 50 -496981
rect -50 -497053 50 -497015
rect -50 -498091 50 -498053
rect -50 -498125 -34 -498091
rect 34 -498125 50 -498091
rect -50 -498141 50 -498125
rect -50 -498199 50 -498183
rect -50 -498233 -34 -498199
rect 34 -498233 50 -498199
rect -50 -498271 50 -498233
rect -50 -499309 50 -499271
rect -50 -499343 -34 -499309
rect 34 -499343 50 -499309
rect -50 -499359 50 -499343
rect -50 -499417 50 -499401
rect -50 -499451 -34 -499417
rect 34 -499451 50 -499417
rect -50 -499489 50 -499451
rect -50 -500527 50 -500489
rect -50 -500561 -34 -500527
rect 34 -500561 50 -500527
rect -50 -500577 50 -500561
rect -50 -500635 50 -500619
rect -50 -500669 -34 -500635
rect 34 -500669 50 -500635
rect -50 -500707 50 -500669
rect -50 -501745 50 -501707
rect -50 -501779 -34 -501745
rect 34 -501779 50 -501745
rect -50 -501795 50 -501779
rect -50 -501853 50 -501837
rect -50 -501887 -34 -501853
rect 34 -501887 50 -501853
rect -50 -501925 50 -501887
rect -50 -502963 50 -502925
rect -50 -502997 -34 -502963
rect 34 -502997 50 -502963
rect -50 -503013 50 -502997
rect -50 -503071 50 -503055
rect -50 -503105 -34 -503071
rect 34 -503105 50 -503071
rect -50 -503143 50 -503105
rect -50 -504181 50 -504143
rect -50 -504215 -34 -504181
rect 34 -504215 50 -504181
rect -50 -504231 50 -504215
rect -50 -504289 50 -504273
rect -50 -504323 -34 -504289
rect 34 -504323 50 -504289
rect -50 -504361 50 -504323
rect -50 -505399 50 -505361
rect -50 -505433 -34 -505399
rect 34 -505433 50 -505399
rect -50 -505449 50 -505433
rect -50 -505507 50 -505491
rect -50 -505541 -34 -505507
rect 34 -505541 50 -505507
rect -50 -505579 50 -505541
rect -50 -506617 50 -506579
rect -50 -506651 -34 -506617
rect 34 -506651 50 -506617
rect -50 -506667 50 -506651
rect -50 -506725 50 -506709
rect -50 -506759 -34 -506725
rect 34 -506759 50 -506725
rect -50 -506797 50 -506759
rect -50 -507835 50 -507797
rect -50 -507869 -34 -507835
rect 34 -507869 50 -507835
rect -50 -507885 50 -507869
rect -50 -507943 50 -507927
rect -50 -507977 -34 -507943
rect 34 -507977 50 -507943
rect -50 -508015 50 -507977
rect -50 -509053 50 -509015
rect -50 -509087 -34 -509053
rect 34 -509087 50 -509053
rect -50 -509103 50 -509087
rect -50 -509161 50 -509145
rect -50 -509195 -34 -509161
rect 34 -509195 50 -509161
rect -50 -509233 50 -509195
rect -50 -510271 50 -510233
rect -50 -510305 -34 -510271
rect 34 -510305 50 -510271
rect -50 -510321 50 -510305
rect -50 -510379 50 -510363
rect -50 -510413 -34 -510379
rect 34 -510413 50 -510379
rect -50 -510451 50 -510413
rect -50 -511489 50 -511451
rect -50 -511523 -34 -511489
rect 34 -511523 50 -511489
rect -50 -511539 50 -511523
rect -50 -511597 50 -511581
rect -50 -511631 -34 -511597
rect 34 -511631 50 -511597
rect -50 -511669 50 -511631
rect -50 -512707 50 -512669
rect -50 -512741 -34 -512707
rect 34 -512741 50 -512707
rect -50 -512757 50 -512741
rect -50 -512815 50 -512799
rect -50 -512849 -34 -512815
rect 34 -512849 50 -512815
rect -50 -512887 50 -512849
rect -50 -513925 50 -513887
rect -50 -513959 -34 -513925
rect 34 -513959 50 -513925
rect -50 -513975 50 -513959
rect -50 -514033 50 -514017
rect -50 -514067 -34 -514033
rect 34 -514067 50 -514033
rect -50 -514105 50 -514067
rect -50 -515143 50 -515105
rect -50 -515177 -34 -515143
rect 34 -515177 50 -515143
rect -50 -515193 50 -515177
rect -50 -515251 50 -515235
rect -50 -515285 -34 -515251
rect 34 -515285 50 -515251
rect -50 -515323 50 -515285
rect -50 -516361 50 -516323
rect -50 -516395 -34 -516361
rect 34 -516395 50 -516361
rect -50 -516411 50 -516395
rect -50 -516469 50 -516453
rect -50 -516503 -34 -516469
rect 34 -516503 50 -516469
rect -50 -516541 50 -516503
rect -50 -517579 50 -517541
rect -50 -517613 -34 -517579
rect 34 -517613 50 -517579
rect -50 -517629 50 -517613
rect -50 -517687 50 -517671
rect -50 -517721 -34 -517687
rect 34 -517721 50 -517687
rect -50 -517759 50 -517721
rect -50 -518797 50 -518759
rect -50 -518831 -34 -518797
rect 34 -518831 50 -518797
rect -50 -518847 50 -518831
rect -50 -518905 50 -518889
rect -50 -518939 -34 -518905
rect 34 -518939 50 -518905
rect -50 -518977 50 -518939
rect -50 -520015 50 -519977
rect -50 -520049 -34 -520015
rect 34 -520049 50 -520015
rect -50 -520065 50 -520049
rect -50 -520123 50 -520107
rect -50 -520157 -34 -520123
rect 34 -520157 50 -520123
rect -50 -520195 50 -520157
rect -50 -521233 50 -521195
rect -50 -521267 -34 -521233
rect 34 -521267 50 -521233
rect -50 -521283 50 -521267
rect -50 -521341 50 -521325
rect -50 -521375 -34 -521341
rect 34 -521375 50 -521341
rect -50 -521413 50 -521375
rect -50 -522451 50 -522413
rect -50 -522485 -34 -522451
rect 34 -522485 50 -522451
rect -50 -522501 50 -522485
rect -50 -522559 50 -522543
rect -50 -522593 -34 -522559
rect 34 -522593 50 -522559
rect -50 -522631 50 -522593
rect -50 -523669 50 -523631
rect -50 -523703 -34 -523669
rect 34 -523703 50 -523669
rect -50 -523719 50 -523703
rect -50 -523777 50 -523761
rect -50 -523811 -34 -523777
rect 34 -523811 50 -523777
rect -50 -523849 50 -523811
rect -50 -524887 50 -524849
rect -50 -524921 -34 -524887
rect 34 -524921 50 -524887
rect -50 -524937 50 -524921
rect -50 -524995 50 -524979
rect -50 -525029 -34 -524995
rect 34 -525029 50 -524995
rect -50 -525067 50 -525029
rect -50 -526105 50 -526067
rect -50 -526139 -34 -526105
rect 34 -526139 50 -526105
rect -50 -526155 50 -526139
rect -50 -526213 50 -526197
rect -50 -526247 -34 -526213
rect 34 -526247 50 -526213
rect -50 -526285 50 -526247
rect -50 -527323 50 -527285
rect -50 -527357 -34 -527323
rect 34 -527357 50 -527323
rect -50 -527373 50 -527357
rect -50 -527431 50 -527415
rect -50 -527465 -34 -527431
rect 34 -527465 50 -527431
rect -50 -527503 50 -527465
rect -50 -528541 50 -528503
rect -50 -528575 -34 -528541
rect 34 -528575 50 -528541
rect -50 -528591 50 -528575
rect -50 -528649 50 -528633
rect -50 -528683 -34 -528649
rect 34 -528683 50 -528649
rect -50 -528721 50 -528683
rect -50 -529759 50 -529721
rect -50 -529793 -34 -529759
rect 34 -529793 50 -529759
rect -50 -529809 50 -529793
rect -50 -529867 50 -529851
rect -50 -529901 -34 -529867
rect 34 -529901 50 -529867
rect -50 -529939 50 -529901
rect -50 -530977 50 -530939
rect -50 -531011 -34 -530977
rect 34 -531011 50 -530977
rect -50 -531027 50 -531011
rect -50 -531085 50 -531069
rect -50 -531119 -34 -531085
rect 34 -531119 50 -531085
rect -50 -531157 50 -531119
rect -50 -532195 50 -532157
rect -50 -532229 -34 -532195
rect 34 -532229 50 -532195
rect -50 -532245 50 -532229
rect -50 -532303 50 -532287
rect -50 -532337 -34 -532303
rect 34 -532337 50 -532303
rect -50 -532375 50 -532337
rect -50 -533413 50 -533375
rect -50 -533447 -34 -533413
rect 34 -533447 50 -533413
rect -50 -533463 50 -533447
rect -50 -533521 50 -533505
rect -50 -533555 -34 -533521
rect 34 -533555 50 -533521
rect -50 -533593 50 -533555
rect -50 -534631 50 -534593
rect -50 -534665 -34 -534631
rect 34 -534665 50 -534631
rect -50 -534681 50 -534665
rect -50 -534739 50 -534723
rect -50 -534773 -34 -534739
rect 34 -534773 50 -534739
rect -50 -534811 50 -534773
rect -50 -535849 50 -535811
rect -50 -535883 -34 -535849
rect 34 -535883 50 -535849
rect -50 -535899 50 -535883
rect -50 -535957 50 -535941
rect -50 -535991 -34 -535957
rect 34 -535991 50 -535957
rect -50 -536029 50 -535991
rect -50 -537067 50 -537029
rect -50 -537101 -34 -537067
rect 34 -537101 50 -537067
rect -50 -537117 50 -537101
rect -50 -537175 50 -537159
rect -50 -537209 -34 -537175
rect 34 -537209 50 -537175
rect -50 -537247 50 -537209
rect -50 -538285 50 -538247
rect -50 -538319 -34 -538285
rect 34 -538319 50 -538285
rect -50 -538335 50 -538319
rect -50 -538393 50 -538377
rect -50 -538427 -34 -538393
rect 34 -538427 50 -538393
rect -50 -538465 50 -538427
rect -50 -539503 50 -539465
rect -50 -539537 -34 -539503
rect 34 -539537 50 -539503
rect -50 -539553 50 -539537
rect -50 -539611 50 -539595
rect -50 -539645 -34 -539611
rect 34 -539645 50 -539611
rect -50 -539683 50 -539645
rect -50 -540721 50 -540683
rect -50 -540755 -34 -540721
rect 34 -540755 50 -540721
rect -50 -540771 50 -540755
rect -50 -540829 50 -540813
rect -50 -540863 -34 -540829
rect 34 -540863 50 -540829
rect -50 -540901 50 -540863
rect -50 -541939 50 -541901
rect -50 -541973 -34 -541939
rect 34 -541973 50 -541939
rect -50 -541989 50 -541973
rect -50 -542047 50 -542031
rect -50 -542081 -34 -542047
rect 34 -542081 50 -542047
rect -50 -542119 50 -542081
rect -50 -543157 50 -543119
rect -50 -543191 -34 -543157
rect 34 -543191 50 -543157
rect -50 -543207 50 -543191
rect -50 -543265 50 -543249
rect -50 -543299 -34 -543265
rect 34 -543299 50 -543265
rect -50 -543337 50 -543299
rect -50 -544375 50 -544337
rect -50 -544409 -34 -544375
rect 34 -544409 50 -544375
rect -50 -544425 50 -544409
rect -50 -544483 50 -544467
rect -50 -544517 -34 -544483
rect 34 -544517 50 -544483
rect -50 -544555 50 -544517
rect -50 -545593 50 -545555
rect -50 -545627 -34 -545593
rect 34 -545627 50 -545593
rect -50 -545643 50 -545627
rect -50 -545701 50 -545685
rect -50 -545735 -34 -545701
rect 34 -545735 50 -545701
rect -50 -545773 50 -545735
rect -50 -546811 50 -546773
rect -50 -546845 -34 -546811
rect 34 -546845 50 -546811
rect -50 -546861 50 -546845
rect -50 -546919 50 -546903
rect -50 -546953 -34 -546919
rect 34 -546953 50 -546919
rect -50 -546991 50 -546953
rect -50 -548029 50 -547991
rect -50 -548063 -34 -548029
rect 34 -548063 50 -548029
rect -50 -548079 50 -548063
rect -50 -548137 50 -548121
rect -50 -548171 -34 -548137
rect 34 -548171 50 -548137
rect -50 -548209 50 -548171
rect -50 -549247 50 -549209
rect -50 -549281 -34 -549247
rect 34 -549281 50 -549247
rect -50 -549297 50 -549281
rect -50 -549355 50 -549339
rect -50 -549389 -34 -549355
rect 34 -549389 50 -549355
rect -50 -549427 50 -549389
rect -50 -550465 50 -550427
rect -50 -550499 -34 -550465
rect 34 -550499 50 -550465
rect -50 -550515 50 -550499
rect -50 -550573 50 -550557
rect -50 -550607 -34 -550573
rect 34 -550607 50 -550573
rect -50 -550645 50 -550607
rect -50 -551683 50 -551645
rect -50 -551717 -34 -551683
rect 34 -551717 50 -551683
rect -50 -551733 50 -551717
rect -50 -551791 50 -551775
rect -50 -551825 -34 -551791
rect 34 -551825 50 -551791
rect -50 -551863 50 -551825
rect -50 -552901 50 -552863
rect -50 -552935 -34 -552901
rect 34 -552935 50 -552901
rect -50 -552951 50 -552935
rect -50 -553009 50 -552993
rect -50 -553043 -34 -553009
rect 34 -553043 50 -553009
rect -50 -553081 50 -553043
rect -50 -554119 50 -554081
rect -50 -554153 -34 -554119
rect 34 -554153 50 -554119
rect -50 -554169 50 -554153
rect -50 -554227 50 -554211
rect -50 -554261 -34 -554227
rect 34 -554261 50 -554227
rect -50 -554299 50 -554261
rect -50 -555337 50 -555299
rect -50 -555371 -34 -555337
rect 34 -555371 50 -555337
rect -50 -555387 50 -555371
rect -50 -555445 50 -555429
rect -50 -555479 -34 -555445
rect 34 -555479 50 -555445
rect -50 -555517 50 -555479
rect -50 -556555 50 -556517
rect -50 -556589 -34 -556555
rect 34 -556589 50 -556555
rect -50 -556605 50 -556589
rect -50 -556663 50 -556647
rect -50 -556697 -34 -556663
rect 34 -556697 50 -556663
rect -50 -556735 50 -556697
rect -50 -557773 50 -557735
rect -50 -557807 -34 -557773
rect 34 -557807 50 -557773
rect -50 -557823 50 -557807
rect -50 -557881 50 -557865
rect -50 -557915 -34 -557881
rect 34 -557915 50 -557881
rect -50 -557953 50 -557915
rect -50 -558991 50 -558953
rect -50 -559025 -34 -558991
rect 34 -559025 50 -558991
rect -50 -559041 50 -559025
rect -50 -559099 50 -559083
rect -50 -559133 -34 -559099
rect 34 -559133 50 -559099
rect -50 -559171 50 -559133
rect -50 -560209 50 -560171
rect -50 -560243 -34 -560209
rect 34 -560243 50 -560209
rect -50 -560259 50 -560243
rect -50 -560317 50 -560301
rect -50 -560351 -34 -560317
rect 34 -560351 50 -560317
rect -50 -560389 50 -560351
rect -50 -561427 50 -561389
rect -50 -561461 -34 -561427
rect 34 -561461 50 -561427
rect -50 -561477 50 -561461
rect -50 -561535 50 -561519
rect -50 -561569 -34 -561535
rect 34 -561569 50 -561535
rect -50 -561607 50 -561569
rect -50 -562645 50 -562607
rect -50 -562679 -34 -562645
rect 34 -562679 50 -562645
rect -50 -562695 50 -562679
rect -50 -562753 50 -562737
rect -50 -562787 -34 -562753
rect 34 -562787 50 -562753
rect -50 -562825 50 -562787
rect -50 -563863 50 -563825
rect -50 -563897 -34 -563863
rect 34 -563897 50 -563863
rect -50 -563913 50 -563897
rect -50 -563971 50 -563955
rect -50 -564005 -34 -563971
rect 34 -564005 50 -563971
rect -50 -564043 50 -564005
rect -50 -565081 50 -565043
rect -50 -565115 -34 -565081
rect 34 -565115 50 -565081
rect -50 -565131 50 -565115
rect -50 -565189 50 -565173
rect -50 -565223 -34 -565189
rect 34 -565223 50 -565189
rect -50 -565261 50 -565223
rect -50 -566299 50 -566261
rect -50 -566333 -34 -566299
rect 34 -566333 50 -566299
rect -50 -566349 50 -566333
rect -50 -566407 50 -566391
rect -50 -566441 -34 -566407
rect 34 -566441 50 -566407
rect -50 -566479 50 -566441
rect -50 -567517 50 -567479
rect -50 -567551 -34 -567517
rect 34 -567551 50 -567517
rect -50 -567567 50 -567551
rect -50 -567625 50 -567609
rect -50 -567659 -34 -567625
rect 34 -567659 50 -567625
rect -50 -567697 50 -567659
rect -50 -568735 50 -568697
rect -50 -568769 -34 -568735
rect 34 -568769 50 -568735
rect -50 -568785 50 -568769
rect -50 -568843 50 -568827
rect -50 -568877 -34 -568843
rect 34 -568877 50 -568843
rect -50 -568915 50 -568877
rect -50 -569953 50 -569915
rect -50 -569987 -34 -569953
rect 34 -569987 50 -569953
rect -50 -570003 50 -569987
rect -50 -570061 50 -570045
rect -50 -570095 -34 -570061
rect 34 -570095 50 -570061
rect -50 -570133 50 -570095
rect -50 -571171 50 -571133
rect -50 -571205 -34 -571171
rect 34 -571205 50 -571171
rect -50 -571221 50 -571205
rect -50 -571279 50 -571263
rect -50 -571313 -34 -571279
rect 34 -571313 50 -571279
rect -50 -571351 50 -571313
rect -50 -572389 50 -572351
rect -50 -572423 -34 -572389
rect 34 -572423 50 -572389
rect -50 -572439 50 -572423
rect -50 -572497 50 -572481
rect -50 -572531 -34 -572497
rect 34 -572531 50 -572497
rect -50 -572569 50 -572531
rect -50 -573607 50 -573569
rect -50 -573641 -34 -573607
rect 34 -573641 50 -573607
rect -50 -573657 50 -573641
rect -50 -573715 50 -573699
rect -50 -573749 -34 -573715
rect 34 -573749 50 -573715
rect -50 -573787 50 -573749
rect -50 -574825 50 -574787
rect -50 -574859 -34 -574825
rect 34 -574859 50 -574825
rect -50 -574875 50 -574859
rect -50 -574933 50 -574917
rect -50 -574967 -34 -574933
rect 34 -574967 50 -574933
rect -50 -575005 50 -574967
rect -50 -576043 50 -576005
rect -50 -576077 -34 -576043
rect 34 -576077 50 -576043
rect -50 -576093 50 -576077
rect -50 -576151 50 -576135
rect -50 -576185 -34 -576151
rect 34 -576185 50 -576151
rect -50 -576223 50 -576185
rect -50 -577261 50 -577223
rect -50 -577295 -34 -577261
rect 34 -577295 50 -577261
rect -50 -577311 50 -577295
rect -50 -577369 50 -577353
rect -50 -577403 -34 -577369
rect 34 -577403 50 -577369
rect -50 -577441 50 -577403
rect -50 -578479 50 -578441
rect -50 -578513 -34 -578479
rect 34 -578513 50 -578479
rect -50 -578529 50 -578513
rect -50 -578587 50 -578571
rect -50 -578621 -34 -578587
rect 34 -578621 50 -578587
rect -50 -578659 50 -578621
rect -50 -579697 50 -579659
rect -50 -579731 -34 -579697
rect 34 -579731 50 -579697
rect -50 -579747 50 -579731
rect -50 -579805 50 -579789
rect -50 -579839 -34 -579805
rect 34 -579839 50 -579805
rect -50 -579877 50 -579839
rect -50 -580915 50 -580877
rect -50 -580949 -34 -580915
rect 34 -580949 50 -580915
rect -50 -580965 50 -580949
rect -50 -581023 50 -581007
rect -50 -581057 -34 -581023
rect 34 -581057 50 -581023
rect -50 -581095 50 -581057
rect -50 -582133 50 -582095
rect -50 -582167 -34 -582133
rect 34 -582167 50 -582133
rect -50 -582183 50 -582167
rect -50 -582241 50 -582225
rect -50 -582275 -34 -582241
rect 34 -582275 50 -582241
rect -50 -582313 50 -582275
rect -50 -583351 50 -583313
rect -50 -583385 -34 -583351
rect 34 -583385 50 -583351
rect -50 -583401 50 -583385
rect -50 -583459 50 -583443
rect -50 -583493 -34 -583459
rect 34 -583493 50 -583459
rect -50 -583531 50 -583493
rect -50 -584569 50 -584531
rect -50 -584603 -34 -584569
rect 34 -584603 50 -584569
rect -50 -584619 50 -584603
rect -50 -584677 50 -584661
rect -50 -584711 -34 -584677
rect 34 -584711 50 -584677
rect -50 -584749 50 -584711
rect -50 -585787 50 -585749
rect -50 -585821 -34 -585787
rect 34 -585821 50 -585787
rect -50 -585837 50 -585821
rect -50 -585895 50 -585879
rect -50 -585929 -34 -585895
rect 34 -585929 50 -585895
rect -50 -585967 50 -585929
rect -50 -587005 50 -586967
rect -50 -587039 -34 -587005
rect 34 -587039 50 -587005
rect -50 -587055 50 -587039
rect -50 -587113 50 -587097
rect -50 -587147 -34 -587113
rect 34 -587147 50 -587113
rect -50 -587185 50 -587147
rect -50 -588223 50 -588185
rect -50 -588257 -34 -588223
rect 34 -588257 50 -588223
rect -50 -588273 50 -588257
rect -50 -588331 50 -588315
rect -50 -588365 -34 -588331
rect 34 -588365 50 -588331
rect -50 -588403 50 -588365
rect -50 -589441 50 -589403
rect -50 -589475 -34 -589441
rect 34 -589475 50 -589441
rect -50 -589491 50 -589475
rect -50 -589549 50 -589533
rect -50 -589583 -34 -589549
rect 34 -589583 50 -589549
rect -50 -589621 50 -589583
rect -50 -590659 50 -590621
rect -50 -590693 -34 -590659
rect 34 -590693 50 -590659
rect -50 -590709 50 -590693
rect -50 -590767 50 -590751
rect -50 -590801 -34 -590767
rect 34 -590801 50 -590767
rect -50 -590839 50 -590801
rect -50 -591877 50 -591839
rect -50 -591911 -34 -591877
rect 34 -591911 50 -591877
rect -50 -591927 50 -591911
rect -50 -591985 50 -591969
rect -50 -592019 -34 -591985
rect 34 -592019 50 -591985
rect -50 -592057 50 -592019
rect -50 -593095 50 -593057
rect -50 -593129 -34 -593095
rect 34 -593129 50 -593095
rect -50 -593145 50 -593129
rect -50 -593203 50 -593187
rect -50 -593237 -34 -593203
rect 34 -593237 50 -593203
rect -50 -593275 50 -593237
rect -50 -594313 50 -594275
rect -50 -594347 -34 -594313
rect 34 -594347 50 -594313
rect -50 -594363 50 -594347
rect -50 -594421 50 -594405
rect -50 -594455 -34 -594421
rect 34 -594455 50 -594421
rect -50 -594493 50 -594455
rect -50 -595531 50 -595493
rect -50 -595565 -34 -595531
rect 34 -595565 50 -595531
rect -50 -595581 50 -595565
rect -50 -595639 50 -595623
rect -50 -595673 -34 -595639
rect 34 -595673 50 -595639
rect -50 -595711 50 -595673
rect -50 -596749 50 -596711
rect -50 -596783 -34 -596749
rect 34 -596783 50 -596749
rect -50 -596799 50 -596783
rect -50 -596857 50 -596841
rect -50 -596891 -34 -596857
rect 34 -596891 50 -596857
rect -50 -596929 50 -596891
rect -50 -597967 50 -597929
rect -50 -598001 -34 -597967
rect 34 -598001 50 -597967
rect -50 -598017 50 -598001
rect -50 -598075 50 -598059
rect -50 -598109 -34 -598075
rect 34 -598109 50 -598075
rect -50 -598147 50 -598109
rect -50 -599185 50 -599147
rect -50 -599219 -34 -599185
rect 34 -599219 50 -599185
rect -50 -599235 50 -599219
rect -50 -599293 50 -599277
rect -50 -599327 -34 -599293
rect 34 -599327 50 -599293
rect -50 -599365 50 -599327
rect -50 -600403 50 -600365
rect -50 -600437 -34 -600403
rect 34 -600437 50 -600403
rect -50 -600453 50 -600437
rect -50 -600511 50 -600495
rect -50 -600545 -34 -600511
rect 34 -600545 50 -600511
rect -50 -600583 50 -600545
rect -50 -601621 50 -601583
rect -50 -601655 -34 -601621
rect 34 -601655 50 -601621
rect -50 -601671 50 -601655
rect -50 -601729 50 -601713
rect -50 -601763 -34 -601729
rect 34 -601763 50 -601729
rect -50 -601801 50 -601763
rect -50 -602839 50 -602801
rect -50 -602873 -34 -602839
rect 34 -602873 50 -602839
rect -50 -602889 50 -602873
rect -50 -602947 50 -602931
rect -50 -602981 -34 -602947
rect 34 -602981 50 -602947
rect -50 -603019 50 -602981
rect -50 -604057 50 -604019
rect -50 -604091 -34 -604057
rect 34 -604091 50 -604057
rect -50 -604107 50 -604091
rect -50 -604165 50 -604149
rect -50 -604199 -34 -604165
rect 34 -604199 50 -604165
rect -50 -604237 50 -604199
rect -50 -605275 50 -605237
rect -50 -605309 -34 -605275
rect 34 -605309 50 -605275
rect -50 -605325 50 -605309
rect -50 -605383 50 -605367
rect -50 -605417 -34 -605383
rect 34 -605417 50 -605383
rect -50 -605455 50 -605417
rect -50 -606493 50 -606455
rect -50 -606527 -34 -606493
rect 34 -606527 50 -606493
rect -50 -606543 50 -606527
rect -50 -606601 50 -606585
rect -50 -606635 -34 -606601
rect 34 -606635 50 -606601
rect -50 -606673 50 -606635
rect -50 -607711 50 -607673
rect -50 -607745 -34 -607711
rect 34 -607745 50 -607711
rect -50 -607761 50 -607745
rect -50 -607819 50 -607803
rect -50 -607853 -34 -607819
rect 34 -607853 50 -607819
rect -50 -607891 50 -607853
rect -50 -608929 50 -608891
rect -50 -608963 -34 -608929
rect 34 -608963 50 -608929
rect -50 -608979 50 -608963
<< polycont >>
rect -34 608929 34 608963
rect -34 607819 34 607853
rect -34 607711 34 607745
rect -34 606601 34 606635
rect -34 606493 34 606527
rect -34 605383 34 605417
rect -34 605275 34 605309
rect -34 604165 34 604199
rect -34 604057 34 604091
rect -34 602947 34 602981
rect -34 602839 34 602873
rect -34 601729 34 601763
rect -34 601621 34 601655
rect -34 600511 34 600545
rect -34 600403 34 600437
rect -34 599293 34 599327
rect -34 599185 34 599219
rect -34 598075 34 598109
rect -34 597967 34 598001
rect -34 596857 34 596891
rect -34 596749 34 596783
rect -34 595639 34 595673
rect -34 595531 34 595565
rect -34 594421 34 594455
rect -34 594313 34 594347
rect -34 593203 34 593237
rect -34 593095 34 593129
rect -34 591985 34 592019
rect -34 591877 34 591911
rect -34 590767 34 590801
rect -34 590659 34 590693
rect -34 589549 34 589583
rect -34 589441 34 589475
rect -34 588331 34 588365
rect -34 588223 34 588257
rect -34 587113 34 587147
rect -34 587005 34 587039
rect -34 585895 34 585929
rect -34 585787 34 585821
rect -34 584677 34 584711
rect -34 584569 34 584603
rect -34 583459 34 583493
rect -34 583351 34 583385
rect -34 582241 34 582275
rect -34 582133 34 582167
rect -34 581023 34 581057
rect -34 580915 34 580949
rect -34 579805 34 579839
rect -34 579697 34 579731
rect -34 578587 34 578621
rect -34 578479 34 578513
rect -34 577369 34 577403
rect -34 577261 34 577295
rect -34 576151 34 576185
rect -34 576043 34 576077
rect -34 574933 34 574967
rect -34 574825 34 574859
rect -34 573715 34 573749
rect -34 573607 34 573641
rect -34 572497 34 572531
rect -34 572389 34 572423
rect -34 571279 34 571313
rect -34 571171 34 571205
rect -34 570061 34 570095
rect -34 569953 34 569987
rect -34 568843 34 568877
rect -34 568735 34 568769
rect -34 567625 34 567659
rect -34 567517 34 567551
rect -34 566407 34 566441
rect -34 566299 34 566333
rect -34 565189 34 565223
rect -34 565081 34 565115
rect -34 563971 34 564005
rect -34 563863 34 563897
rect -34 562753 34 562787
rect -34 562645 34 562679
rect -34 561535 34 561569
rect -34 561427 34 561461
rect -34 560317 34 560351
rect -34 560209 34 560243
rect -34 559099 34 559133
rect -34 558991 34 559025
rect -34 557881 34 557915
rect -34 557773 34 557807
rect -34 556663 34 556697
rect -34 556555 34 556589
rect -34 555445 34 555479
rect -34 555337 34 555371
rect -34 554227 34 554261
rect -34 554119 34 554153
rect -34 553009 34 553043
rect -34 552901 34 552935
rect -34 551791 34 551825
rect -34 551683 34 551717
rect -34 550573 34 550607
rect -34 550465 34 550499
rect -34 549355 34 549389
rect -34 549247 34 549281
rect -34 548137 34 548171
rect -34 548029 34 548063
rect -34 546919 34 546953
rect -34 546811 34 546845
rect -34 545701 34 545735
rect -34 545593 34 545627
rect -34 544483 34 544517
rect -34 544375 34 544409
rect -34 543265 34 543299
rect -34 543157 34 543191
rect -34 542047 34 542081
rect -34 541939 34 541973
rect -34 540829 34 540863
rect -34 540721 34 540755
rect -34 539611 34 539645
rect -34 539503 34 539537
rect -34 538393 34 538427
rect -34 538285 34 538319
rect -34 537175 34 537209
rect -34 537067 34 537101
rect -34 535957 34 535991
rect -34 535849 34 535883
rect -34 534739 34 534773
rect -34 534631 34 534665
rect -34 533521 34 533555
rect -34 533413 34 533447
rect -34 532303 34 532337
rect -34 532195 34 532229
rect -34 531085 34 531119
rect -34 530977 34 531011
rect -34 529867 34 529901
rect -34 529759 34 529793
rect -34 528649 34 528683
rect -34 528541 34 528575
rect -34 527431 34 527465
rect -34 527323 34 527357
rect -34 526213 34 526247
rect -34 526105 34 526139
rect -34 524995 34 525029
rect -34 524887 34 524921
rect -34 523777 34 523811
rect -34 523669 34 523703
rect -34 522559 34 522593
rect -34 522451 34 522485
rect -34 521341 34 521375
rect -34 521233 34 521267
rect -34 520123 34 520157
rect -34 520015 34 520049
rect -34 518905 34 518939
rect -34 518797 34 518831
rect -34 517687 34 517721
rect -34 517579 34 517613
rect -34 516469 34 516503
rect -34 516361 34 516395
rect -34 515251 34 515285
rect -34 515143 34 515177
rect -34 514033 34 514067
rect -34 513925 34 513959
rect -34 512815 34 512849
rect -34 512707 34 512741
rect -34 511597 34 511631
rect -34 511489 34 511523
rect -34 510379 34 510413
rect -34 510271 34 510305
rect -34 509161 34 509195
rect -34 509053 34 509087
rect -34 507943 34 507977
rect -34 507835 34 507869
rect -34 506725 34 506759
rect -34 506617 34 506651
rect -34 505507 34 505541
rect -34 505399 34 505433
rect -34 504289 34 504323
rect -34 504181 34 504215
rect -34 503071 34 503105
rect -34 502963 34 502997
rect -34 501853 34 501887
rect -34 501745 34 501779
rect -34 500635 34 500669
rect -34 500527 34 500561
rect -34 499417 34 499451
rect -34 499309 34 499343
rect -34 498199 34 498233
rect -34 498091 34 498125
rect -34 496981 34 497015
rect -34 496873 34 496907
rect -34 495763 34 495797
rect -34 495655 34 495689
rect -34 494545 34 494579
rect -34 494437 34 494471
rect -34 493327 34 493361
rect -34 493219 34 493253
rect -34 492109 34 492143
rect -34 492001 34 492035
rect -34 490891 34 490925
rect -34 490783 34 490817
rect -34 489673 34 489707
rect -34 489565 34 489599
rect -34 488455 34 488489
rect -34 488347 34 488381
rect -34 487237 34 487271
rect -34 487129 34 487163
rect -34 486019 34 486053
rect -34 485911 34 485945
rect -34 484801 34 484835
rect -34 484693 34 484727
rect -34 483583 34 483617
rect -34 483475 34 483509
rect -34 482365 34 482399
rect -34 482257 34 482291
rect -34 481147 34 481181
rect -34 481039 34 481073
rect -34 479929 34 479963
rect -34 479821 34 479855
rect -34 478711 34 478745
rect -34 478603 34 478637
rect -34 477493 34 477527
rect -34 477385 34 477419
rect -34 476275 34 476309
rect -34 476167 34 476201
rect -34 475057 34 475091
rect -34 474949 34 474983
rect -34 473839 34 473873
rect -34 473731 34 473765
rect -34 472621 34 472655
rect -34 472513 34 472547
rect -34 471403 34 471437
rect -34 471295 34 471329
rect -34 470185 34 470219
rect -34 470077 34 470111
rect -34 468967 34 469001
rect -34 468859 34 468893
rect -34 467749 34 467783
rect -34 467641 34 467675
rect -34 466531 34 466565
rect -34 466423 34 466457
rect -34 465313 34 465347
rect -34 465205 34 465239
rect -34 464095 34 464129
rect -34 463987 34 464021
rect -34 462877 34 462911
rect -34 462769 34 462803
rect -34 461659 34 461693
rect -34 461551 34 461585
rect -34 460441 34 460475
rect -34 460333 34 460367
rect -34 459223 34 459257
rect -34 459115 34 459149
rect -34 458005 34 458039
rect -34 457897 34 457931
rect -34 456787 34 456821
rect -34 456679 34 456713
rect -34 455569 34 455603
rect -34 455461 34 455495
rect -34 454351 34 454385
rect -34 454243 34 454277
rect -34 453133 34 453167
rect -34 453025 34 453059
rect -34 451915 34 451949
rect -34 451807 34 451841
rect -34 450697 34 450731
rect -34 450589 34 450623
rect -34 449479 34 449513
rect -34 449371 34 449405
rect -34 448261 34 448295
rect -34 448153 34 448187
rect -34 447043 34 447077
rect -34 446935 34 446969
rect -34 445825 34 445859
rect -34 445717 34 445751
rect -34 444607 34 444641
rect -34 444499 34 444533
rect -34 443389 34 443423
rect -34 443281 34 443315
rect -34 442171 34 442205
rect -34 442063 34 442097
rect -34 440953 34 440987
rect -34 440845 34 440879
rect -34 439735 34 439769
rect -34 439627 34 439661
rect -34 438517 34 438551
rect -34 438409 34 438443
rect -34 437299 34 437333
rect -34 437191 34 437225
rect -34 436081 34 436115
rect -34 435973 34 436007
rect -34 434863 34 434897
rect -34 434755 34 434789
rect -34 433645 34 433679
rect -34 433537 34 433571
rect -34 432427 34 432461
rect -34 432319 34 432353
rect -34 431209 34 431243
rect -34 431101 34 431135
rect -34 429991 34 430025
rect -34 429883 34 429917
rect -34 428773 34 428807
rect -34 428665 34 428699
rect -34 427555 34 427589
rect -34 427447 34 427481
rect -34 426337 34 426371
rect -34 426229 34 426263
rect -34 425119 34 425153
rect -34 425011 34 425045
rect -34 423901 34 423935
rect -34 423793 34 423827
rect -34 422683 34 422717
rect -34 422575 34 422609
rect -34 421465 34 421499
rect -34 421357 34 421391
rect -34 420247 34 420281
rect -34 420139 34 420173
rect -34 419029 34 419063
rect -34 418921 34 418955
rect -34 417811 34 417845
rect -34 417703 34 417737
rect -34 416593 34 416627
rect -34 416485 34 416519
rect -34 415375 34 415409
rect -34 415267 34 415301
rect -34 414157 34 414191
rect -34 414049 34 414083
rect -34 412939 34 412973
rect -34 412831 34 412865
rect -34 411721 34 411755
rect -34 411613 34 411647
rect -34 410503 34 410537
rect -34 410395 34 410429
rect -34 409285 34 409319
rect -34 409177 34 409211
rect -34 408067 34 408101
rect -34 407959 34 407993
rect -34 406849 34 406883
rect -34 406741 34 406775
rect -34 405631 34 405665
rect -34 405523 34 405557
rect -34 404413 34 404447
rect -34 404305 34 404339
rect -34 403195 34 403229
rect -34 403087 34 403121
rect -34 401977 34 402011
rect -34 401869 34 401903
rect -34 400759 34 400793
rect -34 400651 34 400685
rect -34 399541 34 399575
rect -34 399433 34 399467
rect -34 398323 34 398357
rect -34 398215 34 398249
rect -34 397105 34 397139
rect -34 396997 34 397031
rect -34 395887 34 395921
rect -34 395779 34 395813
rect -34 394669 34 394703
rect -34 394561 34 394595
rect -34 393451 34 393485
rect -34 393343 34 393377
rect -34 392233 34 392267
rect -34 392125 34 392159
rect -34 391015 34 391049
rect -34 390907 34 390941
rect -34 389797 34 389831
rect -34 389689 34 389723
rect -34 388579 34 388613
rect -34 388471 34 388505
rect -34 387361 34 387395
rect -34 387253 34 387287
rect -34 386143 34 386177
rect -34 386035 34 386069
rect -34 384925 34 384959
rect -34 384817 34 384851
rect -34 383707 34 383741
rect -34 383599 34 383633
rect -34 382489 34 382523
rect -34 382381 34 382415
rect -34 381271 34 381305
rect -34 381163 34 381197
rect -34 380053 34 380087
rect -34 379945 34 379979
rect -34 378835 34 378869
rect -34 378727 34 378761
rect -34 377617 34 377651
rect -34 377509 34 377543
rect -34 376399 34 376433
rect -34 376291 34 376325
rect -34 375181 34 375215
rect -34 375073 34 375107
rect -34 373963 34 373997
rect -34 373855 34 373889
rect -34 372745 34 372779
rect -34 372637 34 372671
rect -34 371527 34 371561
rect -34 371419 34 371453
rect -34 370309 34 370343
rect -34 370201 34 370235
rect -34 369091 34 369125
rect -34 368983 34 369017
rect -34 367873 34 367907
rect -34 367765 34 367799
rect -34 366655 34 366689
rect -34 366547 34 366581
rect -34 365437 34 365471
rect -34 365329 34 365363
rect -34 364219 34 364253
rect -34 364111 34 364145
rect -34 363001 34 363035
rect -34 362893 34 362927
rect -34 361783 34 361817
rect -34 361675 34 361709
rect -34 360565 34 360599
rect -34 360457 34 360491
rect -34 359347 34 359381
rect -34 359239 34 359273
rect -34 358129 34 358163
rect -34 358021 34 358055
rect -34 356911 34 356945
rect -34 356803 34 356837
rect -34 355693 34 355727
rect -34 355585 34 355619
rect -34 354475 34 354509
rect -34 354367 34 354401
rect -34 353257 34 353291
rect -34 353149 34 353183
rect -34 352039 34 352073
rect -34 351931 34 351965
rect -34 350821 34 350855
rect -34 350713 34 350747
rect -34 349603 34 349637
rect -34 349495 34 349529
rect -34 348385 34 348419
rect -34 348277 34 348311
rect -34 347167 34 347201
rect -34 347059 34 347093
rect -34 345949 34 345983
rect -34 345841 34 345875
rect -34 344731 34 344765
rect -34 344623 34 344657
rect -34 343513 34 343547
rect -34 343405 34 343439
rect -34 342295 34 342329
rect -34 342187 34 342221
rect -34 341077 34 341111
rect -34 340969 34 341003
rect -34 339859 34 339893
rect -34 339751 34 339785
rect -34 338641 34 338675
rect -34 338533 34 338567
rect -34 337423 34 337457
rect -34 337315 34 337349
rect -34 336205 34 336239
rect -34 336097 34 336131
rect -34 334987 34 335021
rect -34 334879 34 334913
rect -34 333769 34 333803
rect -34 333661 34 333695
rect -34 332551 34 332585
rect -34 332443 34 332477
rect -34 331333 34 331367
rect -34 331225 34 331259
rect -34 330115 34 330149
rect -34 330007 34 330041
rect -34 328897 34 328931
rect -34 328789 34 328823
rect -34 327679 34 327713
rect -34 327571 34 327605
rect -34 326461 34 326495
rect -34 326353 34 326387
rect -34 325243 34 325277
rect -34 325135 34 325169
rect -34 324025 34 324059
rect -34 323917 34 323951
rect -34 322807 34 322841
rect -34 322699 34 322733
rect -34 321589 34 321623
rect -34 321481 34 321515
rect -34 320371 34 320405
rect -34 320263 34 320297
rect -34 319153 34 319187
rect -34 319045 34 319079
rect -34 317935 34 317969
rect -34 317827 34 317861
rect -34 316717 34 316751
rect -34 316609 34 316643
rect -34 315499 34 315533
rect -34 315391 34 315425
rect -34 314281 34 314315
rect -34 314173 34 314207
rect -34 313063 34 313097
rect -34 312955 34 312989
rect -34 311845 34 311879
rect -34 311737 34 311771
rect -34 310627 34 310661
rect -34 310519 34 310553
rect -34 309409 34 309443
rect -34 309301 34 309335
rect -34 308191 34 308225
rect -34 308083 34 308117
rect -34 306973 34 307007
rect -34 306865 34 306899
rect -34 305755 34 305789
rect -34 305647 34 305681
rect -34 304537 34 304571
rect -34 304429 34 304463
rect -34 303319 34 303353
rect -34 303211 34 303245
rect -34 302101 34 302135
rect -34 301993 34 302027
rect -34 300883 34 300917
rect -34 300775 34 300809
rect -34 299665 34 299699
rect -34 299557 34 299591
rect -34 298447 34 298481
rect -34 298339 34 298373
rect -34 297229 34 297263
rect -34 297121 34 297155
rect -34 296011 34 296045
rect -34 295903 34 295937
rect -34 294793 34 294827
rect -34 294685 34 294719
rect -34 293575 34 293609
rect -34 293467 34 293501
rect -34 292357 34 292391
rect -34 292249 34 292283
rect -34 291139 34 291173
rect -34 291031 34 291065
rect -34 289921 34 289955
rect -34 289813 34 289847
rect -34 288703 34 288737
rect -34 288595 34 288629
rect -34 287485 34 287519
rect -34 287377 34 287411
rect -34 286267 34 286301
rect -34 286159 34 286193
rect -34 285049 34 285083
rect -34 284941 34 284975
rect -34 283831 34 283865
rect -34 283723 34 283757
rect -34 282613 34 282647
rect -34 282505 34 282539
rect -34 281395 34 281429
rect -34 281287 34 281321
rect -34 280177 34 280211
rect -34 280069 34 280103
rect -34 278959 34 278993
rect -34 278851 34 278885
rect -34 277741 34 277775
rect -34 277633 34 277667
rect -34 276523 34 276557
rect -34 276415 34 276449
rect -34 275305 34 275339
rect -34 275197 34 275231
rect -34 274087 34 274121
rect -34 273979 34 274013
rect -34 272869 34 272903
rect -34 272761 34 272795
rect -34 271651 34 271685
rect -34 271543 34 271577
rect -34 270433 34 270467
rect -34 270325 34 270359
rect -34 269215 34 269249
rect -34 269107 34 269141
rect -34 267997 34 268031
rect -34 267889 34 267923
rect -34 266779 34 266813
rect -34 266671 34 266705
rect -34 265561 34 265595
rect -34 265453 34 265487
rect -34 264343 34 264377
rect -34 264235 34 264269
rect -34 263125 34 263159
rect -34 263017 34 263051
rect -34 261907 34 261941
rect -34 261799 34 261833
rect -34 260689 34 260723
rect -34 260581 34 260615
rect -34 259471 34 259505
rect -34 259363 34 259397
rect -34 258253 34 258287
rect -34 258145 34 258179
rect -34 257035 34 257069
rect -34 256927 34 256961
rect -34 255817 34 255851
rect -34 255709 34 255743
rect -34 254599 34 254633
rect -34 254491 34 254525
rect -34 253381 34 253415
rect -34 253273 34 253307
rect -34 252163 34 252197
rect -34 252055 34 252089
rect -34 250945 34 250979
rect -34 250837 34 250871
rect -34 249727 34 249761
rect -34 249619 34 249653
rect -34 248509 34 248543
rect -34 248401 34 248435
rect -34 247291 34 247325
rect -34 247183 34 247217
rect -34 246073 34 246107
rect -34 245965 34 245999
rect -34 244855 34 244889
rect -34 244747 34 244781
rect -34 243637 34 243671
rect -34 243529 34 243563
rect -34 242419 34 242453
rect -34 242311 34 242345
rect -34 241201 34 241235
rect -34 241093 34 241127
rect -34 239983 34 240017
rect -34 239875 34 239909
rect -34 238765 34 238799
rect -34 238657 34 238691
rect -34 237547 34 237581
rect -34 237439 34 237473
rect -34 236329 34 236363
rect -34 236221 34 236255
rect -34 235111 34 235145
rect -34 235003 34 235037
rect -34 233893 34 233927
rect -34 233785 34 233819
rect -34 232675 34 232709
rect -34 232567 34 232601
rect -34 231457 34 231491
rect -34 231349 34 231383
rect -34 230239 34 230273
rect -34 230131 34 230165
rect -34 229021 34 229055
rect -34 228913 34 228947
rect -34 227803 34 227837
rect -34 227695 34 227729
rect -34 226585 34 226619
rect -34 226477 34 226511
rect -34 225367 34 225401
rect -34 225259 34 225293
rect -34 224149 34 224183
rect -34 224041 34 224075
rect -34 222931 34 222965
rect -34 222823 34 222857
rect -34 221713 34 221747
rect -34 221605 34 221639
rect -34 220495 34 220529
rect -34 220387 34 220421
rect -34 219277 34 219311
rect -34 219169 34 219203
rect -34 218059 34 218093
rect -34 217951 34 217985
rect -34 216841 34 216875
rect -34 216733 34 216767
rect -34 215623 34 215657
rect -34 215515 34 215549
rect -34 214405 34 214439
rect -34 214297 34 214331
rect -34 213187 34 213221
rect -34 213079 34 213113
rect -34 211969 34 212003
rect -34 211861 34 211895
rect -34 210751 34 210785
rect -34 210643 34 210677
rect -34 209533 34 209567
rect -34 209425 34 209459
rect -34 208315 34 208349
rect -34 208207 34 208241
rect -34 207097 34 207131
rect -34 206989 34 207023
rect -34 205879 34 205913
rect -34 205771 34 205805
rect -34 204661 34 204695
rect -34 204553 34 204587
rect -34 203443 34 203477
rect -34 203335 34 203369
rect -34 202225 34 202259
rect -34 202117 34 202151
rect -34 201007 34 201041
rect -34 200899 34 200933
rect -34 199789 34 199823
rect -34 199681 34 199715
rect -34 198571 34 198605
rect -34 198463 34 198497
rect -34 197353 34 197387
rect -34 197245 34 197279
rect -34 196135 34 196169
rect -34 196027 34 196061
rect -34 194917 34 194951
rect -34 194809 34 194843
rect -34 193699 34 193733
rect -34 193591 34 193625
rect -34 192481 34 192515
rect -34 192373 34 192407
rect -34 191263 34 191297
rect -34 191155 34 191189
rect -34 190045 34 190079
rect -34 189937 34 189971
rect -34 188827 34 188861
rect -34 188719 34 188753
rect -34 187609 34 187643
rect -34 187501 34 187535
rect -34 186391 34 186425
rect -34 186283 34 186317
rect -34 185173 34 185207
rect -34 185065 34 185099
rect -34 183955 34 183989
rect -34 183847 34 183881
rect -34 182737 34 182771
rect -34 182629 34 182663
rect -34 181519 34 181553
rect -34 181411 34 181445
rect -34 180301 34 180335
rect -34 180193 34 180227
rect -34 179083 34 179117
rect -34 178975 34 179009
rect -34 177865 34 177899
rect -34 177757 34 177791
rect -34 176647 34 176681
rect -34 176539 34 176573
rect -34 175429 34 175463
rect -34 175321 34 175355
rect -34 174211 34 174245
rect -34 174103 34 174137
rect -34 172993 34 173027
rect -34 172885 34 172919
rect -34 171775 34 171809
rect -34 171667 34 171701
rect -34 170557 34 170591
rect -34 170449 34 170483
rect -34 169339 34 169373
rect -34 169231 34 169265
rect -34 168121 34 168155
rect -34 168013 34 168047
rect -34 166903 34 166937
rect -34 166795 34 166829
rect -34 165685 34 165719
rect -34 165577 34 165611
rect -34 164467 34 164501
rect -34 164359 34 164393
rect -34 163249 34 163283
rect -34 163141 34 163175
rect -34 162031 34 162065
rect -34 161923 34 161957
rect -34 160813 34 160847
rect -34 160705 34 160739
rect -34 159595 34 159629
rect -34 159487 34 159521
rect -34 158377 34 158411
rect -34 158269 34 158303
rect -34 157159 34 157193
rect -34 157051 34 157085
rect -34 155941 34 155975
rect -34 155833 34 155867
rect -34 154723 34 154757
rect -34 154615 34 154649
rect -34 153505 34 153539
rect -34 153397 34 153431
rect -34 152287 34 152321
rect -34 152179 34 152213
rect -34 151069 34 151103
rect -34 150961 34 150995
rect -34 149851 34 149885
rect -34 149743 34 149777
rect -34 148633 34 148667
rect -34 148525 34 148559
rect -34 147415 34 147449
rect -34 147307 34 147341
rect -34 146197 34 146231
rect -34 146089 34 146123
rect -34 144979 34 145013
rect -34 144871 34 144905
rect -34 143761 34 143795
rect -34 143653 34 143687
rect -34 142543 34 142577
rect -34 142435 34 142469
rect -34 141325 34 141359
rect -34 141217 34 141251
rect -34 140107 34 140141
rect -34 139999 34 140033
rect -34 138889 34 138923
rect -34 138781 34 138815
rect -34 137671 34 137705
rect -34 137563 34 137597
rect -34 136453 34 136487
rect -34 136345 34 136379
rect -34 135235 34 135269
rect -34 135127 34 135161
rect -34 134017 34 134051
rect -34 133909 34 133943
rect -34 132799 34 132833
rect -34 132691 34 132725
rect -34 131581 34 131615
rect -34 131473 34 131507
rect -34 130363 34 130397
rect -34 130255 34 130289
rect -34 129145 34 129179
rect -34 129037 34 129071
rect -34 127927 34 127961
rect -34 127819 34 127853
rect -34 126709 34 126743
rect -34 126601 34 126635
rect -34 125491 34 125525
rect -34 125383 34 125417
rect -34 124273 34 124307
rect -34 124165 34 124199
rect -34 123055 34 123089
rect -34 122947 34 122981
rect -34 121837 34 121871
rect -34 121729 34 121763
rect -34 120619 34 120653
rect -34 120511 34 120545
rect -34 119401 34 119435
rect -34 119293 34 119327
rect -34 118183 34 118217
rect -34 118075 34 118109
rect -34 116965 34 116999
rect -34 116857 34 116891
rect -34 115747 34 115781
rect -34 115639 34 115673
rect -34 114529 34 114563
rect -34 114421 34 114455
rect -34 113311 34 113345
rect -34 113203 34 113237
rect -34 112093 34 112127
rect -34 111985 34 112019
rect -34 110875 34 110909
rect -34 110767 34 110801
rect -34 109657 34 109691
rect -34 109549 34 109583
rect -34 108439 34 108473
rect -34 108331 34 108365
rect -34 107221 34 107255
rect -34 107113 34 107147
rect -34 106003 34 106037
rect -34 105895 34 105929
rect -34 104785 34 104819
rect -34 104677 34 104711
rect -34 103567 34 103601
rect -34 103459 34 103493
rect -34 102349 34 102383
rect -34 102241 34 102275
rect -34 101131 34 101165
rect -34 101023 34 101057
rect -34 99913 34 99947
rect -34 99805 34 99839
rect -34 98695 34 98729
rect -34 98587 34 98621
rect -34 97477 34 97511
rect -34 97369 34 97403
rect -34 96259 34 96293
rect -34 96151 34 96185
rect -34 95041 34 95075
rect -34 94933 34 94967
rect -34 93823 34 93857
rect -34 93715 34 93749
rect -34 92605 34 92639
rect -34 92497 34 92531
rect -34 91387 34 91421
rect -34 91279 34 91313
rect -34 90169 34 90203
rect -34 90061 34 90095
rect -34 88951 34 88985
rect -34 88843 34 88877
rect -34 87733 34 87767
rect -34 87625 34 87659
rect -34 86515 34 86549
rect -34 86407 34 86441
rect -34 85297 34 85331
rect -34 85189 34 85223
rect -34 84079 34 84113
rect -34 83971 34 84005
rect -34 82861 34 82895
rect -34 82753 34 82787
rect -34 81643 34 81677
rect -34 81535 34 81569
rect -34 80425 34 80459
rect -34 80317 34 80351
rect -34 79207 34 79241
rect -34 79099 34 79133
rect -34 77989 34 78023
rect -34 77881 34 77915
rect -34 76771 34 76805
rect -34 76663 34 76697
rect -34 75553 34 75587
rect -34 75445 34 75479
rect -34 74335 34 74369
rect -34 74227 34 74261
rect -34 73117 34 73151
rect -34 73009 34 73043
rect -34 71899 34 71933
rect -34 71791 34 71825
rect -34 70681 34 70715
rect -34 70573 34 70607
rect -34 69463 34 69497
rect -34 69355 34 69389
rect -34 68245 34 68279
rect -34 68137 34 68171
rect -34 67027 34 67061
rect -34 66919 34 66953
rect -34 65809 34 65843
rect -34 65701 34 65735
rect -34 64591 34 64625
rect -34 64483 34 64517
rect -34 63373 34 63407
rect -34 63265 34 63299
rect -34 62155 34 62189
rect -34 62047 34 62081
rect -34 60937 34 60971
rect -34 60829 34 60863
rect -34 59719 34 59753
rect -34 59611 34 59645
rect -34 58501 34 58535
rect -34 58393 34 58427
rect -34 57283 34 57317
rect -34 57175 34 57209
rect -34 56065 34 56099
rect -34 55957 34 55991
rect -34 54847 34 54881
rect -34 54739 34 54773
rect -34 53629 34 53663
rect -34 53521 34 53555
rect -34 52411 34 52445
rect -34 52303 34 52337
rect -34 51193 34 51227
rect -34 51085 34 51119
rect -34 49975 34 50009
rect -34 49867 34 49901
rect -34 48757 34 48791
rect -34 48649 34 48683
rect -34 47539 34 47573
rect -34 47431 34 47465
rect -34 46321 34 46355
rect -34 46213 34 46247
rect -34 45103 34 45137
rect -34 44995 34 45029
rect -34 43885 34 43919
rect -34 43777 34 43811
rect -34 42667 34 42701
rect -34 42559 34 42593
rect -34 41449 34 41483
rect -34 41341 34 41375
rect -34 40231 34 40265
rect -34 40123 34 40157
rect -34 39013 34 39047
rect -34 38905 34 38939
rect -34 37795 34 37829
rect -34 37687 34 37721
rect -34 36577 34 36611
rect -34 36469 34 36503
rect -34 35359 34 35393
rect -34 35251 34 35285
rect -34 34141 34 34175
rect -34 34033 34 34067
rect -34 32923 34 32957
rect -34 32815 34 32849
rect -34 31705 34 31739
rect -34 31597 34 31631
rect -34 30487 34 30521
rect -34 30379 34 30413
rect -34 29269 34 29303
rect -34 29161 34 29195
rect -34 28051 34 28085
rect -34 27943 34 27977
rect -34 26833 34 26867
rect -34 26725 34 26759
rect -34 25615 34 25649
rect -34 25507 34 25541
rect -34 24397 34 24431
rect -34 24289 34 24323
rect -34 23179 34 23213
rect -34 23071 34 23105
rect -34 21961 34 21995
rect -34 21853 34 21887
rect -34 20743 34 20777
rect -34 20635 34 20669
rect -34 19525 34 19559
rect -34 19417 34 19451
rect -34 18307 34 18341
rect -34 18199 34 18233
rect -34 17089 34 17123
rect -34 16981 34 17015
rect -34 15871 34 15905
rect -34 15763 34 15797
rect -34 14653 34 14687
rect -34 14545 34 14579
rect -34 13435 34 13469
rect -34 13327 34 13361
rect -34 12217 34 12251
rect -34 12109 34 12143
rect -34 10999 34 11033
rect -34 10891 34 10925
rect -34 9781 34 9815
rect -34 9673 34 9707
rect -34 8563 34 8597
rect -34 8455 34 8489
rect -34 7345 34 7379
rect -34 7237 34 7271
rect -34 6127 34 6161
rect -34 6019 34 6053
rect -34 4909 34 4943
rect -34 4801 34 4835
rect -34 3691 34 3725
rect -34 3583 34 3617
rect -34 2473 34 2507
rect -34 2365 34 2399
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -34 -2399 34 -2365
rect -34 -2507 34 -2473
rect -34 -3617 34 -3583
rect -34 -3725 34 -3691
rect -34 -4835 34 -4801
rect -34 -4943 34 -4909
rect -34 -6053 34 -6019
rect -34 -6161 34 -6127
rect -34 -7271 34 -7237
rect -34 -7379 34 -7345
rect -34 -8489 34 -8455
rect -34 -8597 34 -8563
rect -34 -9707 34 -9673
rect -34 -9815 34 -9781
rect -34 -10925 34 -10891
rect -34 -11033 34 -10999
rect -34 -12143 34 -12109
rect -34 -12251 34 -12217
rect -34 -13361 34 -13327
rect -34 -13469 34 -13435
rect -34 -14579 34 -14545
rect -34 -14687 34 -14653
rect -34 -15797 34 -15763
rect -34 -15905 34 -15871
rect -34 -17015 34 -16981
rect -34 -17123 34 -17089
rect -34 -18233 34 -18199
rect -34 -18341 34 -18307
rect -34 -19451 34 -19417
rect -34 -19559 34 -19525
rect -34 -20669 34 -20635
rect -34 -20777 34 -20743
rect -34 -21887 34 -21853
rect -34 -21995 34 -21961
rect -34 -23105 34 -23071
rect -34 -23213 34 -23179
rect -34 -24323 34 -24289
rect -34 -24431 34 -24397
rect -34 -25541 34 -25507
rect -34 -25649 34 -25615
rect -34 -26759 34 -26725
rect -34 -26867 34 -26833
rect -34 -27977 34 -27943
rect -34 -28085 34 -28051
rect -34 -29195 34 -29161
rect -34 -29303 34 -29269
rect -34 -30413 34 -30379
rect -34 -30521 34 -30487
rect -34 -31631 34 -31597
rect -34 -31739 34 -31705
rect -34 -32849 34 -32815
rect -34 -32957 34 -32923
rect -34 -34067 34 -34033
rect -34 -34175 34 -34141
rect -34 -35285 34 -35251
rect -34 -35393 34 -35359
rect -34 -36503 34 -36469
rect -34 -36611 34 -36577
rect -34 -37721 34 -37687
rect -34 -37829 34 -37795
rect -34 -38939 34 -38905
rect -34 -39047 34 -39013
rect -34 -40157 34 -40123
rect -34 -40265 34 -40231
rect -34 -41375 34 -41341
rect -34 -41483 34 -41449
rect -34 -42593 34 -42559
rect -34 -42701 34 -42667
rect -34 -43811 34 -43777
rect -34 -43919 34 -43885
rect -34 -45029 34 -44995
rect -34 -45137 34 -45103
rect -34 -46247 34 -46213
rect -34 -46355 34 -46321
rect -34 -47465 34 -47431
rect -34 -47573 34 -47539
rect -34 -48683 34 -48649
rect -34 -48791 34 -48757
rect -34 -49901 34 -49867
rect -34 -50009 34 -49975
rect -34 -51119 34 -51085
rect -34 -51227 34 -51193
rect -34 -52337 34 -52303
rect -34 -52445 34 -52411
rect -34 -53555 34 -53521
rect -34 -53663 34 -53629
rect -34 -54773 34 -54739
rect -34 -54881 34 -54847
rect -34 -55991 34 -55957
rect -34 -56099 34 -56065
rect -34 -57209 34 -57175
rect -34 -57317 34 -57283
rect -34 -58427 34 -58393
rect -34 -58535 34 -58501
rect -34 -59645 34 -59611
rect -34 -59753 34 -59719
rect -34 -60863 34 -60829
rect -34 -60971 34 -60937
rect -34 -62081 34 -62047
rect -34 -62189 34 -62155
rect -34 -63299 34 -63265
rect -34 -63407 34 -63373
rect -34 -64517 34 -64483
rect -34 -64625 34 -64591
rect -34 -65735 34 -65701
rect -34 -65843 34 -65809
rect -34 -66953 34 -66919
rect -34 -67061 34 -67027
rect -34 -68171 34 -68137
rect -34 -68279 34 -68245
rect -34 -69389 34 -69355
rect -34 -69497 34 -69463
rect -34 -70607 34 -70573
rect -34 -70715 34 -70681
rect -34 -71825 34 -71791
rect -34 -71933 34 -71899
rect -34 -73043 34 -73009
rect -34 -73151 34 -73117
rect -34 -74261 34 -74227
rect -34 -74369 34 -74335
rect -34 -75479 34 -75445
rect -34 -75587 34 -75553
rect -34 -76697 34 -76663
rect -34 -76805 34 -76771
rect -34 -77915 34 -77881
rect -34 -78023 34 -77989
rect -34 -79133 34 -79099
rect -34 -79241 34 -79207
rect -34 -80351 34 -80317
rect -34 -80459 34 -80425
rect -34 -81569 34 -81535
rect -34 -81677 34 -81643
rect -34 -82787 34 -82753
rect -34 -82895 34 -82861
rect -34 -84005 34 -83971
rect -34 -84113 34 -84079
rect -34 -85223 34 -85189
rect -34 -85331 34 -85297
rect -34 -86441 34 -86407
rect -34 -86549 34 -86515
rect -34 -87659 34 -87625
rect -34 -87767 34 -87733
rect -34 -88877 34 -88843
rect -34 -88985 34 -88951
rect -34 -90095 34 -90061
rect -34 -90203 34 -90169
rect -34 -91313 34 -91279
rect -34 -91421 34 -91387
rect -34 -92531 34 -92497
rect -34 -92639 34 -92605
rect -34 -93749 34 -93715
rect -34 -93857 34 -93823
rect -34 -94967 34 -94933
rect -34 -95075 34 -95041
rect -34 -96185 34 -96151
rect -34 -96293 34 -96259
rect -34 -97403 34 -97369
rect -34 -97511 34 -97477
rect -34 -98621 34 -98587
rect -34 -98729 34 -98695
rect -34 -99839 34 -99805
rect -34 -99947 34 -99913
rect -34 -101057 34 -101023
rect -34 -101165 34 -101131
rect -34 -102275 34 -102241
rect -34 -102383 34 -102349
rect -34 -103493 34 -103459
rect -34 -103601 34 -103567
rect -34 -104711 34 -104677
rect -34 -104819 34 -104785
rect -34 -105929 34 -105895
rect -34 -106037 34 -106003
rect -34 -107147 34 -107113
rect -34 -107255 34 -107221
rect -34 -108365 34 -108331
rect -34 -108473 34 -108439
rect -34 -109583 34 -109549
rect -34 -109691 34 -109657
rect -34 -110801 34 -110767
rect -34 -110909 34 -110875
rect -34 -112019 34 -111985
rect -34 -112127 34 -112093
rect -34 -113237 34 -113203
rect -34 -113345 34 -113311
rect -34 -114455 34 -114421
rect -34 -114563 34 -114529
rect -34 -115673 34 -115639
rect -34 -115781 34 -115747
rect -34 -116891 34 -116857
rect -34 -116999 34 -116965
rect -34 -118109 34 -118075
rect -34 -118217 34 -118183
rect -34 -119327 34 -119293
rect -34 -119435 34 -119401
rect -34 -120545 34 -120511
rect -34 -120653 34 -120619
rect -34 -121763 34 -121729
rect -34 -121871 34 -121837
rect -34 -122981 34 -122947
rect -34 -123089 34 -123055
rect -34 -124199 34 -124165
rect -34 -124307 34 -124273
rect -34 -125417 34 -125383
rect -34 -125525 34 -125491
rect -34 -126635 34 -126601
rect -34 -126743 34 -126709
rect -34 -127853 34 -127819
rect -34 -127961 34 -127927
rect -34 -129071 34 -129037
rect -34 -129179 34 -129145
rect -34 -130289 34 -130255
rect -34 -130397 34 -130363
rect -34 -131507 34 -131473
rect -34 -131615 34 -131581
rect -34 -132725 34 -132691
rect -34 -132833 34 -132799
rect -34 -133943 34 -133909
rect -34 -134051 34 -134017
rect -34 -135161 34 -135127
rect -34 -135269 34 -135235
rect -34 -136379 34 -136345
rect -34 -136487 34 -136453
rect -34 -137597 34 -137563
rect -34 -137705 34 -137671
rect -34 -138815 34 -138781
rect -34 -138923 34 -138889
rect -34 -140033 34 -139999
rect -34 -140141 34 -140107
rect -34 -141251 34 -141217
rect -34 -141359 34 -141325
rect -34 -142469 34 -142435
rect -34 -142577 34 -142543
rect -34 -143687 34 -143653
rect -34 -143795 34 -143761
rect -34 -144905 34 -144871
rect -34 -145013 34 -144979
rect -34 -146123 34 -146089
rect -34 -146231 34 -146197
rect -34 -147341 34 -147307
rect -34 -147449 34 -147415
rect -34 -148559 34 -148525
rect -34 -148667 34 -148633
rect -34 -149777 34 -149743
rect -34 -149885 34 -149851
rect -34 -150995 34 -150961
rect -34 -151103 34 -151069
rect -34 -152213 34 -152179
rect -34 -152321 34 -152287
rect -34 -153431 34 -153397
rect -34 -153539 34 -153505
rect -34 -154649 34 -154615
rect -34 -154757 34 -154723
rect -34 -155867 34 -155833
rect -34 -155975 34 -155941
rect -34 -157085 34 -157051
rect -34 -157193 34 -157159
rect -34 -158303 34 -158269
rect -34 -158411 34 -158377
rect -34 -159521 34 -159487
rect -34 -159629 34 -159595
rect -34 -160739 34 -160705
rect -34 -160847 34 -160813
rect -34 -161957 34 -161923
rect -34 -162065 34 -162031
rect -34 -163175 34 -163141
rect -34 -163283 34 -163249
rect -34 -164393 34 -164359
rect -34 -164501 34 -164467
rect -34 -165611 34 -165577
rect -34 -165719 34 -165685
rect -34 -166829 34 -166795
rect -34 -166937 34 -166903
rect -34 -168047 34 -168013
rect -34 -168155 34 -168121
rect -34 -169265 34 -169231
rect -34 -169373 34 -169339
rect -34 -170483 34 -170449
rect -34 -170591 34 -170557
rect -34 -171701 34 -171667
rect -34 -171809 34 -171775
rect -34 -172919 34 -172885
rect -34 -173027 34 -172993
rect -34 -174137 34 -174103
rect -34 -174245 34 -174211
rect -34 -175355 34 -175321
rect -34 -175463 34 -175429
rect -34 -176573 34 -176539
rect -34 -176681 34 -176647
rect -34 -177791 34 -177757
rect -34 -177899 34 -177865
rect -34 -179009 34 -178975
rect -34 -179117 34 -179083
rect -34 -180227 34 -180193
rect -34 -180335 34 -180301
rect -34 -181445 34 -181411
rect -34 -181553 34 -181519
rect -34 -182663 34 -182629
rect -34 -182771 34 -182737
rect -34 -183881 34 -183847
rect -34 -183989 34 -183955
rect -34 -185099 34 -185065
rect -34 -185207 34 -185173
rect -34 -186317 34 -186283
rect -34 -186425 34 -186391
rect -34 -187535 34 -187501
rect -34 -187643 34 -187609
rect -34 -188753 34 -188719
rect -34 -188861 34 -188827
rect -34 -189971 34 -189937
rect -34 -190079 34 -190045
rect -34 -191189 34 -191155
rect -34 -191297 34 -191263
rect -34 -192407 34 -192373
rect -34 -192515 34 -192481
rect -34 -193625 34 -193591
rect -34 -193733 34 -193699
rect -34 -194843 34 -194809
rect -34 -194951 34 -194917
rect -34 -196061 34 -196027
rect -34 -196169 34 -196135
rect -34 -197279 34 -197245
rect -34 -197387 34 -197353
rect -34 -198497 34 -198463
rect -34 -198605 34 -198571
rect -34 -199715 34 -199681
rect -34 -199823 34 -199789
rect -34 -200933 34 -200899
rect -34 -201041 34 -201007
rect -34 -202151 34 -202117
rect -34 -202259 34 -202225
rect -34 -203369 34 -203335
rect -34 -203477 34 -203443
rect -34 -204587 34 -204553
rect -34 -204695 34 -204661
rect -34 -205805 34 -205771
rect -34 -205913 34 -205879
rect -34 -207023 34 -206989
rect -34 -207131 34 -207097
rect -34 -208241 34 -208207
rect -34 -208349 34 -208315
rect -34 -209459 34 -209425
rect -34 -209567 34 -209533
rect -34 -210677 34 -210643
rect -34 -210785 34 -210751
rect -34 -211895 34 -211861
rect -34 -212003 34 -211969
rect -34 -213113 34 -213079
rect -34 -213221 34 -213187
rect -34 -214331 34 -214297
rect -34 -214439 34 -214405
rect -34 -215549 34 -215515
rect -34 -215657 34 -215623
rect -34 -216767 34 -216733
rect -34 -216875 34 -216841
rect -34 -217985 34 -217951
rect -34 -218093 34 -218059
rect -34 -219203 34 -219169
rect -34 -219311 34 -219277
rect -34 -220421 34 -220387
rect -34 -220529 34 -220495
rect -34 -221639 34 -221605
rect -34 -221747 34 -221713
rect -34 -222857 34 -222823
rect -34 -222965 34 -222931
rect -34 -224075 34 -224041
rect -34 -224183 34 -224149
rect -34 -225293 34 -225259
rect -34 -225401 34 -225367
rect -34 -226511 34 -226477
rect -34 -226619 34 -226585
rect -34 -227729 34 -227695
rect -34 -227837 34 -227803
rect -34 -228947 34 -228913
rect -34 -229055 34 -229021
rect -34 -230165 34 -230131
rect -34 -230273 34 -230239
rect -34 -231383 34 -231349
rect -34 -231491 34 -231457
rect -34 -232601 34 -232567
rect -34 -232709 34 -232675
rect -34 -233819 34 -233785
rect -34 -233927 34 -233893
rect -34 -235037 34 -235003
rect -34 -235145 34 -235111
rect -34 -236255 34 -236221
rect -34 -236363 34 -236329
rect -34 -237473 34 -237439
rect -34 -237581 34 -237547
rect -34 -238691 34 -238657
rect -34 -238799 34 -238765
rect -34 -239909 34 -239875
rect -34 -240017 34 -239983
rect -34 -241127 34 -241093
rect -34 -241235 34 -241201
rect -34 -242345 34 -242311
rect -34 -242453 34 -242419
rect -34 -243563 34 -243529
rect -34 -243671 34 -243637
rect -34 -244781 34 -244747
rect -34 -244889 34 -244855
rect -34 -245999 34 -245965
rect -34 -246107 34 -246073
rect -34 -247217 34 -247183
rect -34 -247325 34 -247291
rect -34 -248435 34 -248401
rect -34 -248543 34 -248509
rect -34 -249653 34 -249619
rect -34 -249761 34 -249727
rect -34 -250871 34 -250837
rect -34 -250979 34 -250945
rect -34 -252089 34 -252055
rect -34 -252197 34 -252163
rect -34 -253307 34 -253273
rect -34 -253415 34 -253381
rect -34 -254525 34 -254491
rect -34 -254633 34 -254599
rect -34 -255743 34 -255709
rect -34 -255851 34 -255817
rect -34 -256961 34 -256927
rect -34 -257069 34 -257035
rect -34 -258179 34 -258145
rect -34 -258287 34 -258253
rect -34 -259397 34 -259363
rect -34 -259505 34 -259471
rect -34 -260615 34 -260581
rect -34 -260723 34 -260689
rect -34 -261833 34 -261799
rect -34 -261941 34 -261907
rect -34 -263051 34 -263017
rect -34 -263159 34 -263125
rect -34 -264269 34 -264235
rect -34 -264377 34 -264343
rect -34 -265487 34 -265453
rect -34 -265595 34 -265561
rect -34 -266705 34 -266671
rect -34 -266813 34 -266779
rect -34 -267923 34 -267889
rect -34 -268031 34 -267997
rect -34 -269141 34 -269107
rect -34 -269249 34 -269215
rect -34 -270359 34 -270325
rect -34 -270467 34 -270433
rect -34 -271577 34 -271543
rect -34 -271685 34 -271651
rect -34 -272795 34 -272761
rect -34 -272903 34 -272869
rect -34 -274013 34 -273979
rect -34 -274121 34 -274087
rect -34 -275231 34 -275197
rect -34 -275339 34 -275305
rect -34 -276449 34 -276415
rect -34 -276557 34 -276523
rect -34 -277667 34 -277633
rect -34 -277775 34 -277741
rect -34 -278885 34 -278851
rect -34 -278993 34 -278959
rect -34 -280103 34 -280069
rect -34 -280211 34 -280177
rect -34 -281321 34 -281287
rect -34 -281429 34 -281395
rect -34 -282539 34 -282505
rect -34 -282647 34 -282613
rect -34 -283757 34 -283723
rect -34 -283865 34 -283831
rect -34 -284975 34 -284941
rect -34 -285083 34 -285049
rect -34 -286193 34 -286159
rect -34 -286301 34 -286267
rect -34 -287411 34 -287377
rect -34 -287519 34 -287485
rect -34 -288629 34 -288595
rect -34 -288737 34 -288703
rect -34 -289847 34 -289813
rect -34 -289955 34 -289921
rect -34 -291065 34 -291031
rect -34 -291173 34 -291139
rect -34 -292283 34 -292249
rect -34 -292391 34 -292357
rect -34 -293501 34 -293467
rect -34 -293609 34 -293575
rect -34 -294719 34 -294685
rect -34 -294827 34 -294793
rect -34 -295937 34 -295903
rect -34 -296045 34 -296011
rect -34 -297155 34 -297121
rect -34 -297263 34 -297229
rect -34 -298373 34 -298339
rect -34 -298481 34 -298447
rect -34 -299591 34 -299557
rect -34 -299699 34 -299665
rect -34 -300809 34 -300775
rect -34 -300917 34 -300883
rect -34 -302027 34 -301993
rect -34 -302135 34 -302101
rect -34 -303245 34 -303211
rect -34 -303353 34 -303319
rect -34 -304463 34 -304429
rect -34 -304571 34 -304537
rect -34 -305681 34 -305647
rect -34 -305789 34 -305755
rect -34 -306899 34 -306865
rect -34 -307007 34 -306973
rect -34 -308117 34 -308083
rect -34 -308225 34 -308191
rect -34 -309335 34 -309301
rect -34 -309443 34 -309409
rect -34 -310553 34 -310519
rect -34 -310661 34 -310627
rect -34 -311771 34 -311737
rect -34 -311879 34 -311845
rect -34 -312989 34 -312955
rect -34 -313097 34 -313063
rect -34 -314207 34 -314173
rect -34 -314315 34 -314281
rect -34 -315425 34 -315391
rect -34 -315533 34 -315499
rect -34 -316643 34 -316609
rect -34 -316751 34 -316717
rect -34 -317861 34 -317827
rect -34 -317969 34 -317935
rect -34 -319079 34 -319045
rect -34 -319187 34 -319153
rect -34 -320297 34 -320263
rect -34 -320405 34 -320371
rect -34 -321515 34 -321481
rect -34 -321623 34 -321589
rect -34 -322733 34 -322699
rect -34 -322841 34 -322807
rect -34 -323951 34 -323917
rect -34 -324059 34 -324025
rect -34 -325169 34 -325135
rect -34 -325277 34 -325243
rect -34 -326387 34 -326353
rect -34 -326495 34 -326461
rect -34 -327605 34 -327571
rect -34 -327713 34 -327679
rect -34 -328823 34 -328789
rect -34 -328931 34 -328897
rect -34 -330041 34 -330007
rect -34 -330149 34 -330115
rect -34 -331259 34 -331225
rect -34 -331367 34 -331333
rect -34 -332477 34 -332443
rect -34 -332585 34 -332551
rect -34 -333695 34 -333661
rect -34 -333803 34 -333769
rect -34 -334913 34 -334879
rect -34 -335021 34 -334987
rect -34 -336131 34 -336097
rect -34 -336239 34 -336205
rect -34 -337349 34 -337315
rect -34 -337457 34 -337423
rect -34 -338567 34 -338533
rect -34 -338675 34 -338641
rect -34 -339785 34 -339751
rect -34 -339893 34 -339859
rect -34 -341003 34 -340969
rect -34 -341111 34 -341077
rect -34 -342221 34 -342187
rect -34 -342329 34 -342295
rect -34 -343439 34 -343405
rect -34 -343547 34 -343513
rect -34 -344657 34 -344623
rect -34 -344765 34 -344731
rect -34 -345875 34 -345841
rect -34 -345983 34 -345949
rect -34 -347093 34 -347059
rect -34 -347201 34 -347167
rect -34 -348311 34 -348277
rect -34 -348419 34 -348385
rect -34 -349529 34 -349495
rect -34 -349637 34 -349603
rect -34 -350747 34 -350713
rect -34 -350855 34 -350821
rect -34 -351965 34 -351931
rect -34 -352073 34 -352039
rect -34 -353183 34 -353149
rect -34 -353291 34 -353257
rect -34 -354401 34 -354367
rect -34 -354509 34 -354475
rect -34 -355619 34 -355585
rect -34 -355727 34 -355693
rect -34 -356837 34 -356803
rect -34 -356945 34 -356911
rect -34 -358055 34 -358021
rect -34 -358163 34 -358129
rect -34 -359273 34 -359239
rect -34 -359381 34 -359347
rect -34 -360491 34 -360457
rect -34 -360599 34 -360565
rect -34 -361709 34 -361675
rect -34 -361817 34 -361783
rect -34 -362927 34 -362893
rect -34 -363035 34 -363001
rect -34 -364145 34 -364111
rect -34 -364253 34 -364219
rect -34 -365363 34 -365329
rect -34 -365471 34 -365437
rect -34 -366581 34 -366547
rect -34 -366689 34 -366655
rect -34 -367799 34 -367765
rect -34 -367907 34 -367873
rect -34 -369017 34 -368983
rect -34 -369125 34 -369091
rect -34 -370235 34 -370201
rect -34 -370343 34 -370309
rect -34 -371453 34 -371419
rect -34 -371561 34 -371527
rect -34 -372671 34 -372637
rect -34 -372779 34 -372745
rect -34 -373889 34 -373855
rect -34 -373997 34 -373963
rect -34 -375107 34 -375073
rect -34 -375215 34 -375181
rect -34 -376325 34 -376291
rect -34 -376433 34 -376399
rect -34 -377543 34 -377509
rect -34 -377651 34 -377617
rect -34 -378761 34 -378727
rect -34 -378869 34 -378835
rect -34 -379979 34 -379945
rect -34 -380087 34 -380053
rect -34 -381197 34 -381163
rect -34 -381305 34 -381271
rect -34 -382415 34 -382381
rect -34 -382523 34 -382489
rect -34 -383633 34 -383599
rect -34 -383741 34 -383707
rect -34 -384851 34 -384817
rect -34 -384959 34 -384925
rect -34 -386069 34 -386035
rect -34 -386177 34 -386143
rect -34 -387287 34 -387253
rect -34 -387395 34 -387361
rect -34 -388505 34 -388471
rect -34 -388613 34 -388579
rect -34 -389723 34 -389689
rect -34 -389831 34 -389797
rect -34 -390941 34 -390907
rect -34 -391049 34 -391015
rect -34 -392159 34 -392125
rect -34 -392267 34 -392233
rect -34 -393377 34 -393343
rect -34 -393485 34 -393451
rect -34 -394595 34 -394561
rect -34 -394703 34 -394669
rect -34 -395813 34 -395779
rect -34 -395921 34 -395887
rect -34 -397031 34 -396997
rect -34 -397139 34 -397105
rect -34 -398249 34 -398215
rect -34 -398357 34 -398323
rect -34 -399467 34 -399433
rect -34 -399575 34 -399541
rect -34 -400685 34 -400651
rect -34 -400793 34 -400759
rect -34 -401903 34 -401869
rect -34 -402011 34 -401977
rect -34 -403121 34 -403087
rect -34 -403229 34 -403195
rect -34 -404339 34 -404305
rect -34 -404447 34 -404413
rect -34 -405557 34 -405523
rect -34 -405665 34 -405631
rect -34 -406775 34 -406741
rect -34 -406883 34 -406849
rect -34 -407993 34 -407959
rect -34 -408101 34 -408067
rect -34 -409211 34 -409177
rect -34 -409319 34 -409285
rect -34 -410429 34 -410395
rect -34 -410537 34 -410503
rect -34 -411647 34 -411613
rect -34 -411755 34 -411721
rect -34 -412865 34 -412831
rect -34 -412973 34 -412939
rect -34 -414083 34 -414049
rect -34 -414191 34 -414157
rect -34 -415301 34 -415267
rect -34 -415409 34 -415375
rect -34 -416519 34 -416485
rect -34 -416627 34 -416593
rect -34 -417737 34 -417703
rect -34 -417845 34 -417811
rect -34 -418955 34 -418921
rect -34 -419063 34 -419029
rect -34 -420173 34 -420139
rect -34 -420281 34 -420247
rect -34 -421391 34 -421357
rect -34 -421499 34 -421465
rect -34 -422609 34 -422575
rect -34 -422717 34 -422683
rect -34 -423827 34 -423793
rect -34 -423935 34 -423901
rect -34 -425045 34 -425011
rect -34 -425153 34 -425119
rect -34 -426263 34 -426229
rect -34 -426371 34 -426337
rect -34 -427481 34 -427447
rect -34 -427589 34 -427555
rect -34 -428699 34 -428665
rect -34 -428807 34 -428773
rect -34 -429917 34 -429883
rect -34 -430025 34 -429991
rect -34 -431135 34 -431101
rect -34 -431243 34 -431209
rect -34 -432353 34 -432319
rect -34 -432461 34 -432427
rect -34 -433571 34 -433537
rect -34 -433679 34 -433645
rect -34 -434789 34 -434755
rect -34 -434897 34 -434863
rect -34 -436007 34 -435973
rect -34 -436115 34 -436081
rect -34 -437225 34 -437191
rect -34 -437333 34 -437299
rect -34 -438443 34 -438409
rect -34 -438551 34 -438517
rect -34 -439661 34 -439627
rect -34 -439769 34 -439735
rect -34 -440879 34 -440845
rect -34 -440987 34 -440953
rect -34 -442097 34 -442063
rect -34 -442205 34 -442171
rect -34 -443315 34 -443281
rect -34 -443423 34 -443389
rect -34 -444533 34 -444499
rect -34 -444641 34 -444607
rect -34 -445751 34 -445717
rect -34 -445859 34 -445825
rect -34 -446969 34 -446935
rect -34 -447077 34 -447043
rect -34 -448187 34 -448153
rect -34 -448295 34 -448261
rect -34 -449405 34 -449371
rect -34 -449513 34 -449479
rect -34 -450623 34 -450589
rect -34 -450731 34 -450697
rect -34 -451841 34 -451807
rect -34 -451949 34 -451915
rect -34 -453059 34 -453025
rect -34 -453167 34 -453133
rect -34 -454277 34 -454243
rect -34 -454385 34 -454351
rect -34 -455495 34 -455461
rect -34 -455603 34 -455569
rect -34 -456713 34 -456679
rect -34 -456821 34 -456787
rect -34 -457931 34 -457897
rect -34 -458039 34 -458005
rect -34 -459149 34 -459115
rect -34 -459257 34 -459223
rect -34 -460367 34 -460333
rect -34 -460475 34 -460441
rect -34 -461585 34 -461551
rect -34 -461693 34 -461659
rect -34 -462803 34 -462769
rect -34 -462911 34 -462877
rect -34 -464021 34 -463987
rect -34 -464129 34 -464095
rect -34 -465239 34 -465205
rect -34 -465347 34 -465313
rect -34 -466457 34 -466423
rect -34 -466565 34 -466531
rect -34 -467675 34 -467641
rect -34 -467783 34 -467749
rect -34 -468893 34 -468859
rect -34 -469001 34 -468967
rect -34 -470111 34 -470077
rect -34 -470219 34 -470185
rect -34 -471329 34 -471295
rect -34 -471437 34 -471403
rect -34 -472547 34 -472513
rect -34 -472655 34 -472621
rect -34 -473765 34 -473731
rect -34 -473873 34 -473839
rect -34 -474983 34 -474949
rect -34 -475091 34 -475057
rect -34 -476201 34 -476167
rect -34 -476309 34 -476275
rect -34 -477419 34 -477385
rect -34 -477527 34 -477493
rect -34 -478637 34 -478603
rect -34 -478745 34 -478711
rect -34 -479855 34 -479821
rect -34 -479963 34 -479929
rect -34 -481073 34 -481039
rect -34 -481181 34 -481147
rect -34 -482291 34 -482257
rect -34 -482399 34 -482365
rect -34 -483509 34 -483475
rect -34 -483617 34 -483583
rect -34 -484727 34 -484693
rect -34 -484835 34 -484801
rect -34 -485945 34 -485911
rect -34 -486053 34 -486019
rect -34 -487163 34 -487129
rect -34 -487271 34 -487237
rect -34 -488381 34 -488347
rect -34 -488489 34 -488455
rect -34 -489599 34 -489565
rect -34 -489707 34 -489673
rect -34 -490817 34 -490783
rect -34 -490925 34 -490891
rect -34 -492035 34 -492001
rect -34 -492143 34 -492109
rect -34 -493253 34 -493219
rect -34 -493361 34 -493327
rect -34 -494471 34 -494437
rect -34 -494579 34 -494545
rect -34 -495689 34 -495655
rect -34 -495797 34 -495763
rect -34 -496907 34 -496873
rect -34 -497015 34 -496981
rect -34 -498125 34 -498091
rect -34 -498233 34 -498199
rect -34 -499343 34 -499309
rect -34 -499451 34 -499417
rect -34 -500561 34 -500527
rect -34 -500669 34 -500635
rect -34 -501779 34 -501745
rect -34 -501887 34 -501853
rect -34 -502997 34 -502963
rect -34 -503105 34 -503071
rect -34 -504215 34 -504181
rect -34 -504323 34 -504289
rect -34 -505433 34 -505399
rect -34 -505541 34 -505507
rect -34 -506651 34 -506617
rect -34 -506759 34 -506725
rect -34 -507869 34 -507835
rect -34 -507977 34 -507943
rect -34 -509087 34 -509053
rect -34 -509195 34 -509161
rect -34 -510305 34 -510271
rect -34 -510413 34 -510379
rect -34 -511523 34 -511489
rect -34 -511631 34 -511597
rect -34 -512741 34 -512707
rect -34 -512849 34 -512815
rect -34 -513959 34 -513925
rect -34 -514067 34 -514033
rect -34 -515177 34 -515143
rect -34 -515285 34 -515251
rect -34 -516395 34 -516361
rect -34 -516503 34 -516469
rect -34 -517613 34 -517579
rect -34 -517721 34 -517687
rect -34 -518831 34 -518797
rect -34 -518939 34 -518905
rect -34 -520049 34 -520015
rect -34 -520157 34 -520123
rect -34 -521267 34 -521233
rect -34 -521375 34 -521341
rect -34 -522485 34 -522451
rect -34 -522593 34 -522559
rect -34 -523703 34 -523669
rect -34 -523811 34 -523777
rect -34 -524921 34 -524887
rect -34 -525029 34 -524995
rect -34 -526139 34 -526105
rect -34 -526247 34 -526213
rect -34 -527357 34 -527323
rect -34 -527465 34 -527431
rect -34 -528575 34 -528541
rect -34 -528683 34 -528649
rect -34 -529793 34 -529759
rect -34 -529901 34 -529867
rect -34 -531011 34 -530977
rect -34 -531119 34 -531085
rect -34 -532229 34 -532195
rect -34 -532337 34 -532303
rect -34 -533447 34 -533413
rect -34 -533555 34 -533521
rect -34 -534665 34 -534631
rect -34 -534773 34 -534739
rect -34 -535883 34 -535849
rect -34 -535991 34 -535957
rect -34 -537101 34 -537067
rect -34 -537209 34 -537175
rect -34 -538319 34 -538285
rect -34 -538427 34 -538393
rect -34 -539537 34 -539503
rect -34 -539645 34 -539611
rect -34 -540755 34 -540721
rect -34 -540863 34 -540829
rect -34 -541973 34 -541939
rect -34 -542081 34 -542047
rect -34 -543191 34 -543157
rect -34 -543299 34 -543265
rect -34 -544409 34 -544375
rect -34 -544517 34 -544483
rect -34 -545627 34 -545593
rect -34 -545735 34 -545701
rect -34 -546845 34 -546811
rect -34 -546953 34 -546919
rect -34 -548063 34 -548029
rect -34 -548171 34 -548137
rect -34 -549281 34 -549247
rect -34 -549389 34 -549355
rect -34 -550499 34 -550465
rect -34 -550607 34 -550573
rect -34 -551717 34 -551683
rect -34 -551825 34 -551791
rect -34 -552935 34 -552901
rect -34 -553043 34 -553009
rect -34 -554153 34 -554119
rect -34 -554261 34 -554227
rect -34 -555371 34 -555337
rect -34 -555479 34 -555445
rect -34 -556589 34 -556555
rect -34 -556697 34 -556663
rect -34 -557807 34 -557773
rect -34 -557915 34 -557881
rect -34 -559025 34 -558991
rect -34 -559133 34 -559099
rect -34 -560243 34 -560209
rect -34 -560351 34 -560317
rect -34 -561461 34 -561427
rect -34 -561569 34 -561535
rect -34 -562679 34 -562645
rect -34 -562787 34 -562753
rect -34 -563897 34 -563863
rect -34 -564005 34 -563971
rect -34 -565115 34 -565081
rect -34 -565223 34 -565189
rect -34 -566333 34 -566299
rect -34 -566441 34 -566407
rect -34 -567551 34 -567517
rect -34 -567659 34 -567625
rect -34 -568769 34 -568735
rect -34 -568877 34 -568843
rect -34 -569987 34 -569953
rect -34 -570095 34 -570061
rect -34 -571205 34 -571171
rect -34 -571313 34 -571279
rect -34 -572423 34 -572389
rect -34 -572531 34 -572497
rect -34 -573641 34 -573607
rect -34 -573749 34 -573715
rect -34 -574859 34 -574825
rect -34 -574967 34 -574933
rect -34 -576077 34 -576043
rect -34 -576185 34 -576151
rect -34 -577295 34 -577261
rect -34 -577403 34 -577369
rect -34 -578513 34 -578479
rect -34 -578621 34 -578587
rect -34 -579731 34 -579697
rect -34 -579839 34 -579805
rect -34 -580949 34 -580915
rect -34 -581057 34 -581023
rect -34 -582167 34 -582133
rect -34 -582275 34 -582241
rect -34 -583385 34 -583351
rect -34 -583493 34 -583459
rect -34 -584603 34 -584569
rect -34 -584711 34 -584677
rect -34 -585821 34 -585787
rect -34 -585929 34 -585895
rect -34 -587039 34 -587005
rect -34 -587147 34 -587113
rect -34 -588257 34 -588223
rect -34 -588365 34 -588331
rect -34 -589475 34 -589441
rect -34 -589583 34 -589549
rect -34 -590693 34 -590659
rect -34 -590801 34 -590767
rect -34 -591911 34 -591877
rect -34 -592019 34 -591985
rect -34 -593129 34 -593095
rect -34 -593237 34 -593203
rect -34 -594347 34 -594313
rect -34 -594455 34 -594421
rect -34 -595565 34 -595531
rect -34 -595673 34 -595639
rect -34 -596783 34 -596749
rect -34 -596891 34 -596857
rect -34 -598001 34 -597967
rect -34 -598109 34 -598075
rect -34 -599219 34 -599185
rect -34 -599327 34 -599293
rect -34 -600437 34 -600403
rect -34 -600545 34 -600511
rect -34 -601655 34 -601621
rect -34 -601763 34 -601729
rect -34 -602873 34 -602839
rect -34 -602981 34 -602947
rect -34 -604091 34 -604057
rect -34 -604199 34 -604165
rect -34 -605309 34 -605275
rect -34 -605417 34 -605383
rect -34 -606527 34 -606493
rect -34 -606635 34 -606601
rect -34 -607745 34 -607711
rect -34 -607853 34 -607819
rect -34 -608963 34 -608929
<< locali >>
rect -230 609067 -134 609101
rect 134 609067 230 609101
rect -230 609005 -196 609067
rect 196 609005 230 609067
rect -50 608929 -34 608963
rect 34 608929 50 608963
rect -96 608879 -62 608895
rect -96 607887 -62 607903
rect 62 608879 96 608895
rect 62 607887 96 607903
rect -50 607819 -34 607853
rect 34 607819 50 607853
rect -50 607711 -34 607745
rect 34 607711 50 607745
rect -96 607661 -62 607677
rect -96 606669 -62 606685
rect 62 607661 96 607677
rect 62 606669 96 606685
rect -50 606601 -34 606635
rect 34 606601 50 606635
rect -50 606493 -34 606527
rect 34 606493 50 606527
rect -96 606443 -62 606459
rect -96 605451 -62 605467
rect 62 606443 96 606459
rect 62 605451 96 605467
rect -50 605383 -34 605417
rect 34 605383 50 605417
rect -50 605275 -34 605309
rect 34 605275 50 605309
rect -96 605225 -62 605241
rect -96 604233 -62 604249
rect 62 605225 96 605241
rect 62 604233 96 604249
rect -50 604165 -34 604199
rect 34 604165 50 604199
rect -50 604057 -34 604091
rect 34 604057 50 604091
rect -96 604007 -62 604023
rect -96 603015 -62 603031
rect 62 604007 96 604023
rect 62 603015 96 603031
rect -50 602947 -34 602981
rect 34 602947 50 602981
rect -50 602839 -34 602873
rect 34 602839 50 602873
rect -96 602789 -62 602805
rect -96 601797 -62 601813
rect 62 602789 96 602805
rect 62 601797 96 601813
rect -50 601729 -34 601763
rect 34 601729 50 601763
rect -50 601621 -34 601655
rect 34 601621 50 601655
rect -96 601571 -62 601587
rect -96 600579 -62 600595
rect 62 601571 96 601587
rect 62 600579 96 600595
rect -50 600511 -34 600545
rect 34 600511 50 600545
rect -50 600403 -34 600437
rect 34 600403 50 600437
rect -96 600353 -62 600369
rect -96 599361 -62 599377
rect 62 600353 96 600369
rect 62 599361 96 599377
rect -50 599293 -34 599327
rect 34 599293 50 599327
rect -50 599185 -34 599219
rect 34 599185 50 599219
rect -96 599135 -62 599151
rect -96 598143 -62 598159
rect 62 599135 96 599151
rect 62 598143 96 598159
rect -50 598075 -34 598109
rect 34 598075 50 598109
rect -50 597967 -34 598001
rect 34 597967 50 598001
rect -96 597917 -62 597933
rect -96 596925 -62 596941
rect 62 597917 96 597933
rect 62 596925 96 596941
rect -50 596857 -34 596891
rect 34 596857 50 596891
rect -50 596749 -34 596783
rect 34 596749 50 596783
rect -96 596699 -62 596715
rect -96 595707 -62 595723
rect 62 596699 96 596715
rect 62 595707 96 595723
rect -50 595639 -34 595673
rect 34 595639 50 595673
rect -50 595531 -34 595565
rect 34 595531 50 595565
rect -96 595481 -62 595497
rect -96 594489 -62 594505
rect 62 595481 96 595497
rect 62 594489 96 594505
rect -50 594421 -34 594455
rect 34 594421 50 594455
rect -50 594313 -34 594347
rect 34 594313 50 594347
rect -96 594263 -62 594279
rect -96 593271 -62 593287
rect 62 594263 96 594279
rect 62 593271 96 593287
rect -50 593203 -34 593237
rect 34 593203 50 593237
rect -50 593095 -34 593129
rect 34 593095 50 593129
rect -96 593045 -62 593061
rect -96 592053 -62 592069
rect 62 593045 96 593061
rect 62 592053 96 592069
rect -50 591985 -34 592019
rect 34 591985 50 592019
rect -50 591877 -34 591911
rect 34 591877 50 591911
rect -96 591827 -62 591843
rect -96 590835 -62 590851
rect 62 591827 96 591843
rect 62 590835 96 590851
rect -50 590767 -34 590801
rect 34 590767 50 590801
rect -50 590659 -34 590693
rect 34 590659 50 590693
rect -96 590609 -62 590625
rect -96 589617 -62 589633
rect 62 590609 96 590625
rect 62 589617 96 589633
rect -50 589549 -34 589583
rect 34 589549 50 589583
rect -50 589441 -34 589475
rect 34 589441 50 589475
rect -96 589391 -62 589407
rect -96 588399 -62 588415
rect 62 589391 96 589407
rect 62 588399 96 588415
rect -50 588331 -34 588365
rect 34 588331 50 588365
rect -50 588223 -34 588257
rect 34 588223 50 588257
rect -96 588173 -62 588189
rect -96 587181 -62 587197
rect 62 588173 96 588189
rect 62 587181 96 587197
rect -50 587113 -34 587147
rect 34 587113 50 587147
rect -50 587005 -34 587039
rect 34 587005 50 587039
rect -96 586955 -62 586971
rect -96 585963 -62 585979
rect 62 586955 96 586971
rect 62 585963 96 585979
rect -50 585895 -34 585929
rect 34 585895 50 585929
rect -50 585787 -34 585821
rect 34 585787 50 585821
rect -96 585737 -62 585753
rect -96 584745 -62 584761
rect 62 585737 96 585753
rect 62 584745 96 584761
rect -50 584677 -34 584711
rect 34 584677 50 584711
rect -50 584569 -34 584603
rect 34 584569 50 584603
rect -96 584519 -62 584535
rect -96 583527 -62 583543
rect 62 584519 96 584535
rect 62 583527 96 583543
rect -50 583459 -34 583493
rect 34 583459 50 583493
rect -50 583351 -34 583385
rect 34 583351 50 583385
rect -96 583301 -62 583317
rect -96 582309 -62 582325
rect 62 583301 96 583317
rect 62 582309 96 582325
rect -50 582241 -34 582275
rect 34 582241 50 582275
rect -50 582133 -34 582167
rect 34 582133 50 582167
rect -96 582083 -62 582099
rect -96 581091 -62 581107
rect 62 582083 96 582099
rect 62 581091 96 581107
rect -50 581023 -34 581057
rect 34 581023 50 581057
rect -50 580915 -34 580949
rect 34 580915 50 580949
rect -96 580865 -62 580881
rect -96 579873 -62 579889
rect 62 580865 96 580881
rect 62 579873 96 579889
rect -50 579805 -34 579839
rect 34 579805 50 579839
rect -50 579697 -34 579731
rect 34 579697 50 579731
rect -96 579647 -62 579663
rect -96 578655 -62 578671
rect 62 579647 96 579663
rect 62 578655 96 578671
rect -50 578587 -34 578621
rect 34 578587 50 578621
rect -50 578479 -34 578513
rect 34 578479 50 578513
rect -96 578429 -62 578445
rect -96 577437 -62 577453
rect 62 578429 96 578445
rect 62 577437 96 577453
rect -50 577369 -34 577403
rect 34 577369 50 577403
rect -50 577261 -34 577295
rect 34 577261 50 577295
rect -96 577211 -62 577227
rect -96 576219 -62 576235
rect 62 577211 96 577227
rect 62 576219 96 576235
rect -50 576151 -34 576185
rect 34 576151 50 576185
rect -50 576043 -34 576077
rect 34 576043 50 576077
rect -96 575993 -62 576009
rect -96 575001 -62 575017
rect 62 575993 96 576009
rect 62 575001 96 575017
rect -50 574933 -34 574967
rect 34 574933 50 574967
rect -50 574825 -34 574859
rect 34 574825 50 574859
rect -96 574775 -62 574791
rect -96 573783 -62 573799
rect 62 574775 96 574791
rect 62 573783 96 573799
rect -50 573715 -34 573749
rect 34 573715 50 573749
rect -50 573607 -34 573641
rect 34 573607 50 573641
rect -96 573557 -62 573573
rect -96 572565 -62 572581
rect 62 573557 96 573573
rect 62 572565 96 572581
rect -50 572497 -34 572531
rect 34 572497 50 572531
rect -50 572389 -34 572423
rect 34 572389 50 572423
rect -96 572339 -62 572355
rect -96 571347 -62 571363
rect 62 572339 96 572355
rect 62 571347 96 571363
rect -50 571279 -34 571313
rect 34 571279 50 571313
rect -50 571171 -34 571205
rect 34 571171 50 571205
rect -96 571121 -62 571137
rect -96 570129 -62 570145
rect 62 571121 96 571137
rect 62 570129 96 570145
rect -50 570061 -34 570095
rect 34 570061 50 570095
rect -50 569953 -34 569987
rect 34 569953 50 569987
rect -96 569903 -62 569919
rect -96 568911 -62 568927
rect 62 569903 96 569919
rect 62 568911 96 568927
rect -50 568843 -34 568877
rect 34 568843 50 568877
rect -50 568735 -34 568769
rect 34 568735 50 568769
rect -96 568685 -62 568701
rect -96 567693 -62 567709
rect 62 568685 96 568701
rect 62 567693 96 567709
rect -50 567625 -34 567659
rect 34 567625 50 567659
rect -50 567517 -34 567551
rect 34 567517 50 567551
rect -96 567467 -62 567483
rect -96 566475 -62 566491
rect 62 567467 96 567483
rect 62 566475 96 566491
rect -50 566407 -34 566441
rect 34 566407 50 566441
rect -50 566299 -34 566333
rect 34 566299 50 566333
rect -96 566249 -62 566265
rect -96 565257 -62 565273
rect 62 566249 96 566265
rect 62 565257 96 565273
rect -50 565189 -34 565223
rect 34 565189 50 565223
rect -50 565081 -34 565115
rect 34 565081 50 565115
rect -96 565031 -62 565047
rect -96 564039 -62 564055
rect 62 565031 96 565047
rect 62 564039 96 564055
rect -50 563971 -34 564005
rect 34 563971 50 564005
rect -50 563863 -34 563897
rect 34 563863 50 563897
rect -96 563813 -62 563829
rect -96 562821 -62 562837
rect 62 563813 96 563829
rect 62 562821 96 562837
rect -50 562753 -34 562787
rect 34 562753 50 562787
rect -50 562645 -34 562679
rect 34 562645 50 562679
rect -96 562595 -62 562611
rect -96 561603 -62 561619
rect 62 562595 96 562611
rect 62 561603 96 561619
rect -50 561535 -34 561569
rect 34 561535 50 561569
rect -50 561427 -34 561461
rect 34 561427 50 561461
rect -96 561377 -62 561393
rect -96 560385 -62 560401
rect 62 561377 96 561393
rect 62 560385 96 560401
rect -50 560317 -34 560351
rect 34 560317 50 560351
rect -50 560209 -34 560243
rect 34 560209 50 560243
rect -96 560159 -62 560175
rect -96 559167 -62 559183
rect 62 560159 96 560175
rect 62 559167 96 559183
rect -50 559099 -34 559133
rect 34 559099 50 559133
rect -50 558991 -34 559025
rect 34 558991 50 559025
rect -96 558941 -62 558957
rect -96 557949 -62 557965
rect 62 558941 96 558957
rect 62 557949 96 557965
rect -50 557881 -34 557915
rect 34 557881 50 557915
rect -50 557773 -34 557807
rect 34 557773 50 557807
rect -96 557723 -62 557739
rect -96 556731 -62 556747
rect 62 557723 96 557739
rect 62 556731 96 556747
rect -50 556663 -34 556697
rect 34 556663 50 556697
rect -50 556555 -34 556589
rect 34 556555 50 556589
rect -96 556505 -62 556521
rect -96 555513 -62 555529
rect 62 556505 96 556521
rect 62 555513 96 555529
rect -50 555445 -34 555479
rect 34 555445 50 555479
rect -50 555337 -34 555371
rect 34 555337 50 555371
rect -96 555287 -62 555303
rect -96 554295 -62 554311
rect 62 555287 96 555303
rect 62 554295 96 554311
rect -50 554227 -34 554261
rect 34 554227 50 554261
rect -50 554119 -34 554153
rect 34 554119 50 554153
rect -96 554069 -62 554085
rect -96 553077 -62 553093
rect 62 554069 96 554085
rect 62 553077 96 553093
rect -50 553009 -34 553043
rect 34 553009 50 553043
rect -50 552901 -34 552935
rect 34 552901 50 552935
rect -96 552851 -62 552867
rect -96 551859 -62 551875
rect 62 552851 96 552867
rect 62 551859 96 551875
rect -50 551791 -34 551825
rect 34 551791 50 551825
rect -50 551683 -34 551717
rect 34 551683 50 551717
rect -96 551633 -62 551649
rect -96 550641 -62 550657
rect 62 551633 96 551649
rect 62 550641 96 550657
rect -50 550573 -34 550607
rect 34 550573 50 550607
rect -50 550465 -34 550499
rect 34 550465 50 550499
rect -96 550415 -62 550431
rect -96 549423 -62 549439
rect 62 550415 96 550431
rect 62 549423 96 549439
rect -50 549355 -34 549389
rect 34 549355 50 549389
rect -50 549247 -34 549281
rect 34 549247 50 549281
rect -96 549197 -62 549213
rect -96 548205 -62 548221
rect 62 549197 96 549213
rect 62 548205 96 548221
rect -50 548137 -34 548171
rect 34 548137 50 548171
rect -50 548029 -34 548063
rect 34 548029 50 548063
rect -96 547979 -62 547995
rect -96 546987 -62 547003
rect 62 547979 96 547995
rect 62 546987 96 547003
rect -50 546919 -34 546953
rect 34 546919 50 546953
rect -50 546811 -34 546845
rect 34 546811 50 546845
rect -96 546761 -62 546777
rect -96 545769 -62 545785
rect 62 546761 96 546777
rect 62 545769 96 545785
rect -50 545701 -34 545735
rect 34 545701 50 545735
rect -50 545593 -34 545627
rect 34 545593 50 545627
rect -96 545543 -62 545559
rect -96 544551 -62 544567
rect 62 545543 96 545559
rect 62 544551 96 544567
rect -50 544483 -34 544517
rect 34 544483 50 544517
rect -50 544375 -34 544409
rect 34 544375 50 544409
rect -96 544325 -62 544341
rect -96 543333 -62 543349
rect 62 544325 96 544341
rect 62 543333 96 543349
rect -50 543265 -34 543299
rect 34 543265 50 543299
rect -50 543157 -34 543191
rect 34 543157 50 543191
rect -96 543107 -62 543123
rect -96 542115 -62 542131
rect 62 543107 96 543123
rect 62 542115 96 542131
rect -50 542047 -34 542081
rect 34 542047 50 542081
rect -50 541939 -34 541973
rect 34 541939 50 541973
rect -96 541889 -62 541905
rect -96 540897 -62 540913
rect 62 541889 96 541905
rect 62 540897 96 540913
rect -50 540829 -34 540863
rect 34 540829 50 540863
rect -50 540721 -34 540755
rect 34 540721 50 540755
rect -96 540671 -62 540687
rect -96 539679 -62 539695
rect 62 540671 96 540687
rect 62 539679 96 539695
rect -50 539611 -34 539645
rect 34 539611 50 539645
rect -50 539503 -34 539537
rect 34 539503 50 539537
rect -96 539453 -62 539469
rect -96 538461 -62 538477
rect 62 539453 96 539469
rect 62 538461 96 538477
rect -50 538393 -34 538427
rect 34 538393 50 538427
rect -50 538285 -34 538319
rect 34 538285 50 538319
rect -96 538235 -62 538251
rect -96 537243 -62 537259
rect 62 538235 96 538251
rect 62 537243 96 537259
rect -50 537175 -34 537209
rect 34 537175 50 537209
rect -50 537067 -34 537101
rect 34 537067 50 537101
rect -96 537017 -62 537033
rect -96 536025 -62 536041
rect 62 537017 96 537033
rect 62 536025 96 536041
rect -50 535957 -34 535991
rect 34 535957 50 535991
rect -50 535849 -34 535883
rect 34 535849 50 535883
rect -96 535799 -62 535815
rect -96 534807 -62 534823
rect 62 535799 96 535815
rect 62 534807 96 534823
rect -50 534739 -34 534773
rect 34 534739 50 534773
rect -50 534631 -34 534665
rect 34 534631 50 534665
rect -96 534581 -62 534597
rect -96 533589 -62 533605
rect 62 534581 96 534597
rect 62 533589 96 533605
rect -50 533521 -34 533555
rect 34 533521 50 533555
rect -50 533413 -34 533447
rect 34 533413 50 533447
rect -96 533363 -62 533379
rect -96 532371 -62 532387
rect 62 533363 96 533379
rect 62 532371 96 532387
rect -50 532303 -34 532337
rect 34 532303 50 532337
rect -50 532195 -34 532229
rect 34 532195 50 532229
rect -96 532145 -62 532161
rect -96 531153 -62 531169
rect 62 532145 96 532161
rect 62 531153 96 531169
rect -50 531085 -34 531119
rect 34 531085 50 531119
rect -50 530977 -34 531011
rect 34 530977 50 531011
rect -96 530927 -62 530943
rect -96 529935 -62 529951
rect 62 530927 96 530943
rect 62 529935 96 529951
rect -50 529867 -34 529901
rect 34 529867 50 529901
rect -50 529759 -34 529793
rect 34 529759 50 529793
rect -96 529709 -62 529725
rect -96 528717 -62 528733
rect 62 529709 96 529725
rect 62 528717 96 528733
rect -50 528649 -34 528683
rect 34 528649 50 528683
rect -50 528541 -34 528575
rect 34 528541 50 528575
rect -96 528491 -62 528507
rect -96 527499 -62 527515
rect 62 528491 96 528507
rect 62 527499 96 527515
rect -50 527431 -34 527465
rect 34 527431 50 527465
rect -50 527323 -34 527357
rect 34 527323 50 527357
rect -96 527273 -62 527289
rect -96 526281 -62 526297
rect 62 527273 96 527289
rect 62 526281 96 526297
rect -50 526213 -34 526247
rect 34 526213 50 526247
rect -50 526105 -34 526139
rect 34 526105 50 526139
rect -96 526055 -62 526071
rect -96 525063 -62 525079
rect 62 526055 96 526071
rect 62 525063 96 525079
rect -50 524995 -34 525029
rect 34 524995 50 525029
rect -50 524887 -34 524921
rect 34 524887 50 524921
rect -96 524837 -62 524853
rect -96 523845 -62 523861
rect 62 524837 96 524853
rect 62 523845 96 523861
rect -50 523777 -34 523811
rect 34 523777 50 523811
rect -50 523669 -34 523703
rect 34 523669 50 523703
rect -96 523619 -62 523635
rect -96 522627 -62 522643
rect 62 523619 96 523635
rect 62 522627 96 522643
rect -50 522559 -34 522593
rect 34 522559 50 522593
rect -50 522451 -34 522485
rect 34 522451 50 522485
rect -96 522401 -62 522417
rect -96 521409 -62 521425
rect 62 522401 96 522417
rect 62 521409 96 521425
rect -50 521341 -34 521375
rect 34 521341 50 521375
rect -50 521233 -34 521267
rect 34 521233 50 521267
rect -96 521183 -62 521199
rect -96 520191 -62 520207
rect 62 521183 96 521199
rect 62 520191 96 520207
rect -50 520123 -34 520157
rect 34 520123 50 520157
rect -50 520015 -34 520049
rect 34 520015 50 520049
rect -96 519965 -62 519981
rect -96 518973 -62 518989
rect 62 519965 96 519981
rect 62 518973 96 518989
rect -50 518905 -34 518939
rect 34 518905 50 518939
rect -50 518797 -34 518831
rect 34 518797 50 518831
rect -96 518747 -62 518763
rect -96 517755 -62 517771
rect 62 518747 96 518763
rect 62 517755 96 517771
rect -50 517687 -34 517721
rect 34 517687 50 517721
rect -50 517579 -34 517613
rect 34 517579 50 517613
rect -96 517529 -62 517545
rect -96 516537 -62 516553
rect 62 517529 96 517545
rect 62 516537 96 516553
rect -50 516469 -34 516503
rect 34 516469 50 516503
rect -50 516361 -34 516395
rect 34 516361 50 516395
rect -96 516311 -62 516327
rect -96 515319 -62 515335
rect 62 516311 96 516327
rect 62 515319 96 515335
rect -50 515251 -34 515285
rect 34 515251 50 515285
rect -50 515143 -34 515177
rect 34 515143 50 515177
rect -96 515093 -62 515109
rect -96 514101 -62 514117
rect 62 515093 96 515109
rect 62 514101 96 514117
rect -50 514033 -34 514067
rect 34 514033 50 514067
rect -50 513925 -34 513959
rect 34 513925 50 513959
rect -96 513875 -62 513891
rect -96 512883 -62 512899
rect 62 513875 96 513891
rect 62 512883 96 512899
rect -50 512815 -34 512849
rect 34 512815 50 512849
rect -50 512707 -34 512741
rect 34 512707 50 512741
rect -96 512657 -62 512673
rect -96 511665 -62 511681
rect 62 512657 96 512673
rect 62 511665 96 511681
rect -50 511597 -34 511631
rect 34 511597 50 511631
rect -50 511489 -34 511523
rect 34 511489 50 511523
rect -96 511439 -62 511455
rect -96 510447 -62 510463
rect 62 511439 96 511455
rect 62 510447 96 510463
rect -50 510379 -34 510413
rect 34 510379 50 510413
rect -50 510271 -34 510305
rect 34 510271 50 510305
rect -96 510221 -62 510237
rect -96 509229 -62 509245
rect 62 510221 96 510237
rect 62 509229 96 509245
rect -50 509161 -34 509195
rect 34 509161 50 509195
rect -50 509053 -34 509087
rect 34 509053 50 509087
rect -96 509003 -62 509019
rect -96 508011 -62 508027
rect 62 509003 96 509019
rect 62 508011 96 508027
rect -50 507943 -34 507977
rect 34 507943 50 507977
rect -50 507835 -34 507869
rect 34 507835 50 507869
rect -96 507785 -62 507801
rect -96 506793 -62 506809
rect 62 507785 96 507801
rect 62 506793 96 506809
rect -50 506725 -34 506759
rect 34 506725 50 506759
rect -50 506617 -34 506651
rect 34 506617 50 506651
rect -96 506567 -62 506583
rect -96 505575 -62 505591
rect 62 506567 96 506583
rect 62 505575 96 505591
rect -50 505507 -34 505541
rect 34 505507 50 505541
rect -50 505399 -34 505433
rect 34 505399 50 505433
rect -96 505349 -62 505365
rect -96 504357 -62 504373
rect 62 505349 96 505365
rect 62 504357 96 504373
rect -50 504289 -34 504323
rect 34 504289 50 504323
rect -50 504181 -34 504215
rect 34 504181 50 504215
rect -96 504131 -62 504147
rect -96 503139 -62 503155
rect 62 504131 96 504147
rect 62 503139 96 503155
rect -50 503071 -34 503105
rect 34 503071 50 503105
rect -50 502963 -34 502997
rect 34 502963 50 502997
rect -96 502913 -62 502929
rect -96 501921 -62 501937
rect 62 502913 96 502929
rect 62 501921 96 501937
rect -50 501853 -34 501887
rect 34 501853 50 501887
rect -50 501745 -34 501779
rect 34 501745 50 501779
rect -96 501695 -62 501711
rect -96 500703 -62 500719
rect 62 501695 96 501711
rect 62 500703 96 500719
rect -50 500635 -34 500669
rect 34 500635 50 500669
rect -50 500527 -34 500561
rect 34 500527 50 500561
rect -96 500477 -62 500493
rect -96 499485 -62 499501
rect 62 500477 96 500493
rect 62 499485 96 499501
rect -50 499417 -34 499451
rect 34 499417 50 499451
rect -50 499309 -34 499343
rect 34 499309 50 499343
rect -96 499259 -62 499275
rect -96 498267 -62 498283
rect 62 499259 96 499275
rect 62 498267 96 498283
rect -50 498199 -34 498233
rect 34 498199 50 498233
rect -50 498091 -34 498125
rect 34 498091 50 498125
rect -96 498041 -62 498057
rect -96 497049 -62 497065
rect 62 498041 96 498057
rect 62 497049 96 497065
rect -50 496981 -34 497015
rect 34 496981 50 497015
rect -50 496873 -34 496907
rect 34 496873 50 496907
rect -96 496823 -62 496839
rect -96 495831 -62 495847
rect 62 496823 96 496839
rect 62 495831 96 495847
rect -50 495763 -34 495797
rect 34 495763 50 495797
rect -50 495655 -34 495689
rect 34 495655 50 495689
rect -96 495605 -62 495621
rect -96 494613 -62 494629
rect 62 495605 96 495621
rect 62 494613 96 494629
rect -50 494545 -34 494579
rect 34 494545 50 494579
rect -50 494437 -34 494471
rect 34 494437 50 494471
rect -96 494387 -62 494403
rect -96 493395 -62 493411
rect 62 494387 96 494403
rect 62 493395 96 493411
rect -50 493327 -34 493361
rect 34 493327 50 493361
rect -50 493219 -34 493253
rect 34 493219 50 493253
rect -96 493169 -62 493185
rect -96 492177 -62 492193
rect 62 493169 96 493185
rect 62 492177 96 492193
rect -50 492109 -34 492143
rect 34 492109 50 492143
rect -50 492001 -34 492035
rect 34 492001 50 492035
rect -96 491951 -62 491967
rect -96 490959 -62 490975
rect 62 491951 96 491967
rect 62 490959 96 490975
rect -50 490891 -34 490925
rect 34 490891 50 490925
rect -50 490783 -34 490817
rect 34 490783 50 490817
rect -96 490733 -62 490749
rect -96 489741 -62 489757
rect 62 490733 96 490749
rect 62 489741 96 489757
rect -50 489673 -34 489707
rect 34 489673 50 489707
rect -50 489565 -34 489599
rect 34 489565 50 489599
rect -96 489515 -62 489531
rect -96 488523 -62 488539
rect 62 489515 96 489531
rect 62 488523 96 488539
rect -50 488455 -34 488489
rect 34 488455 50 488489
rect -50 488347 -34 488381
rect 34 488347 50 488381
rect -96 488297 -62 488313
rect -96 487305 -62 487321
rect 62 488297 96 488313
rect 62 487305 96 487321
rect -50 487237 -34 487271
rect 34 487237 50 487271
rect -50 487129 -34 487163
rect 34 487129 50 487163
rect -96 487079 -62 487095
rect -96 486087 -62 486103
rect 62 487079 96 487095
rect 62 486087 96 486103
rect -50 486019 -34 486053
rect 34 486019 50 486053
rect -50 485911 -34 485945
rect 34 485911 50 485945
rect -96 485861 -62 485877
rect -96 484869 -62 484885
rect 62 485861 96 485877
rect 62 484869 96 484885
rect -50 484801 -34 484835
rect 34 484801 50 484835
rect -50 484693 -34 484727
rect 34 484693 50 484727
rect -96 484643 -62 484659
rect -96 483651 -62 483667
rect 62 484643 96 484659
rect 62 483651 96 483667
rect -50 483583 -34 483617
rect 34 483583 50 483617
rect -50 483475 -34 483509
rect 34 483475 50 483509
rect -96 483425 -62 483441
rect -96 482433 -62 482449
rect 62 483425 96 483441
rect 62 482433 96 482449
rect -50 482365 -34 482399
rect 34 482365 50 482399
rect -50 482257 -34 482291
rect 34 482257 50 482291
rect -96 482207 -62 482223
rect -96 481215 -62 481231
rect 62 482207 96 482223
rect 62 481215 96 481231
rect -50 481147 -34 481181
rect 34 481147 50 481181
rect -50 481039 -34 481073
rect 34 481039 50 481073
rect -96 480989 -62 481005
rect -96 479997 -62 480013
rect 62 480989 96 481005
rect 62 479997 96 480013
rect -50 479929 -34 479963
rect 34 479929 50 479963
rect -50 479821 -34 479855
rect 34 479821 50 479855
rect -96 479771 -62 479787
rect -96 478779 -62 478795
rect 62 479771 96 479787
rect 62 478779 96 478795
rect -50 478711 -34 478745
rect 34 478711 50 478745
rect -50 478603 -34 478637
rect 34 478603 50 478637
rect -96 478553 -62 478569
rect -96 477561 -62 477577
rect 62 478553 96 478569
rect 62 477561 96 477577
rect -50 477493 -34 477527
rect 34 477493 50 477527
rect -50 477385 -34 477419
rect 34 477385 50 477419
rect -96 477335 -62 477351
rect -96 476343 -62 476359
rect 62 477335 96 477351
rect 62 476343 96 476359
rect -50 476275 -34 476309
rect 34 476275 50 476309
rect -50 476167 -34 476201
rect 34 476167 50 476201
rect -96 476117 -62 476133
rect -96 475125 -62 475141
rect 62 476117 96 476133
rect 62 475125 96 475141
rect -50 475057 -34 475091
rect 34 475057 50 475091
rect -50 474949 -34 474983
rect 34 474949 50 474983
rect -96 474899 -62 474915
rect -96 473907 -62 473923
rect 62 474899 96 474915
rect 62 473907 96 473923
rect -50 473839 -34 473873
rect 34 473839 50 473873
rect -50 473731 -34 473765
rect 34 473731 50 473765
rect -96 473681 -62 473697
rect -96 472689 -62 472705
rect 62 473681 96 473697
rect 62 472689 96 472705
rect -50 472621 -34 472655
rect 34 472621 50 472655
rect -50 472513 -34 472547
rect 34 472513 50 472547
rect -96 472463 -62 472479
rect -96 471471 -62 471487
rect 62 472463 96 472479
rect 62 471471 96 471487
rect -50 471403 -34 471437
rect 34 471403 50 471437
rect -50 471295 -34 471329
rect 34 471295 50 471329
rect -96 471245 -62 471261
rect -96 470253 -62 470269
rect 62 471245 96 471261
rect 62 470253 96 470269
rect -50 470185 -34 470219
rect 34 470185 50 470219
rect -50 470077 -34 470111
rect 34 470077 50 470111
rect -96 470027 -62 470043
rect -96 469035 -62 469051
rect 62 470027 96 470043
rect 62 469035 96 469051
rect -50 468967 -34 469001
rect 34 468967 50 469001
rect -50 468859 -34 468893
rect 34 468859 50 468893
rect -96 468809 -62 468825
rect -96 467817 -62 467833
rect 62 468809 96 468825
rect 62 467817 96 467833
rect -50 467749 -34 467783
rect 34 467749 50 467783
rect -50 467641 -34 467675
rect 34 467641 50 467675
rect -96 467591 -62 467607
rect -96 466599 -62 466615
rect 62 467591 96 467607
rect 62 466599 96 466615
rect -50 466531 -34 466565
rect 34 466531 50 466565
rect -50 466423 -34 466457
rect 34 466423 50 466457
rect -96 466373 -62 466389
rect -96 465381 -62 465397
rect 62 466373 96 466389
rect 62 465381 96 465397
rect -50 465313 -34 465347
rect 34 465313 50 465347
rect -50 465205 -34 465239
rect 34 465205 50 465239
rect -96 465155 -62 465171
rect -96 464163 -62 464179
rect 62 465155 96 465171
rect 62 464163 96 464179
rect -50 464095 -34 464129
rect 34 464095 50 464129
rect -50 463987 -34 464021
rect 34 463987 50 464021
rect -96 463937 -62 463953
rect -96 462945 -62 462961
rect 62 463937 96 463953
rect 62 462945 96 462961
rect -50 462877 -34 462911
rect 34 462877 50 462911
rect -50 462769 -34 462803
rect 34 462769 50 462803
rect -96 462719 -62 462735
rect -96 461727 -62 461743
rect 62 462719 96 462735
rect 62 461727 96 461743
rect -50 461659 -34 461693
rect 34 461659 50 461693
rect -50 461551 -34 461585
rect 34 461551 50 461585
rect -96 461501 -62 461517
rect -96 460509 -62 460525
rect 62 461501 96 461517
rect 62 460509 96 460525
rect -50 460441 -34 460475
rect 34 460441 50 460475
rect -50 460333 -34 460367
rect 34 460333 50 460367
rect -96 460283 -62 460299
rect -96 459291 -62 459307
rect 62 460283 96 460299
rect 62 459291 96 459307
rect -50 459223 -34 459257
rect 34 459223 50 459257
rect -50 459115 -34 459149
rect 34 459115 50 459149
rect -96 459065 -62 459081
rect -96 458073 -62 458089
rect 62 459065 96 459081
rect 62 458073 96 458089
rect -50 458005 -34 458039
rect 34 458005 50 458039
rect -50 457897 -34 457931
rect 34 457897 50 457931
rect -96 457847 -62 457863
rect -96 456855 -62 456871
rect 62 457847 96 457863
rect 62 456855 96 456871
rect -50 456787 -34 456821
rect 34 456787 50 456821
rect -50 456679 -34 456713
rect 34 456679 50 456713
rect -96 456629 -62 456645
rect -96 455637 -62 455653
rect 62 456629 96 456645
rect 62 455637 96 455653
rect -50 455569 -34 455603
rect 34 455569 50 455603
rect -50 455461 -34 455495
rect 34 455461 50 455495
rect -96 455411 -62 455427
rect -96 454419 -62 454435
rect 62 455411 96 455427
rect 62 454419 96 454435
rect -50 454351 -34 454385
rect 34 454351 50 454385
rect -50 454243 -34 454277
rect 34 454243 50 454277
rect -96 454193 -62 454209
rect -96 453201 -62 453217
rect 62 454193 96 454209
rect 62 453201 96 453217
rect -50 453133 -34 453167
rect 34 453133 50 453167
rect -50 453025 -34 453059
rect 34 453025 50 453059
rect -96 452975 -62 452991
rect -96 451983 -62 451999
rect 62 452975 96 452991
rect 62 451983 96 451999
rect -50 451915 -34 451949
rect 34 451915 50 451949
rect -50 451807 -34 451841
rect 34 451807 50 451841
rect -96 451757 -62 451773
rect -96 450765 -62 450781
rect 62 451757 96 451773
rect 62 450765 96 450781
rect -50 450697 -34 450731
rect 34 450697 50 450731
rect -50 450589 -34 450623
rect 34 450589 50 450623
rect -96 450539 -62 450555
rect -96 449547 -62 449563
rect 62 450539 96 450555
rect 62 449547 96 449563
rect -50 449479 -34 449513
rect 34 449479 50 449513
rect -50 449371 -34 449405
rect 34 449371 50 449405
rect -96 449321 -62 449337
rect -96 448329 -62 448345
rect 62 449321 96 449337
rect 62 448329 96 448345
rect -50 448261 -34 448295
rect 34 448261 50 448295
rect -50 448153 -34 448187
rect 34 448153 50 448187
rect -96 448103 -62 448119
rect -96 447111 -62 447127
rect 62 448103 96 448119
rect 62 447111 96 447127
rect -50 447043 -34 447077
rect 34 447043 50 447077
rect -50 446935 -34 446969
rect 34 446935 50 446969
rect -96 446885 -62 446901
rect -96 445893 -62 445909
rect 62 446885 96 446901
rect 62 445893 96 445909
rect -50 445825 -34 445859
rect 34 445825 50 445859
rect -50 445717 -34 445751
rect 34 445717 50 445751
rect -96 445667 -62 445683
rect -96 444675 -62 444691
rect 62 445667 96 445683
rect 62 444675 96 444691
rect -50 444607 -34 444641
rect 34 444607 50 444641
rect -50 444499 -34 444533
rect 34 444499 50 444533
rect -96 444449 -62 444465
rect -96 443457 -62 443473
rect 62 444449 96 444465
rect 62 443457 96 443473
rect -50 443389 -34 443423
rect 34 443389 50 443423
rect -50 443281 -34 443315
rect 34 443281 50 443315
rect -96 443231 -62 443247
rect -96 442239 -62 442255
rect 62 443231 96 443247
rect 62 442239 96 442255
rect -50 442171 -34 442205
rect 34 442171 50 442205
rect -50 442063 -34 442097
rect 34 442063 50 442097
rect -96 442013 -62 442029
rect -96 441021 -62 441037
rect 62 442013 96 442029
rect 62 441021 96 441037
rect -50 440953 -34 440987
rect 34 440953 50 440987
rect -50 440845 -34 440879
rect 34 440845 50 440879
rect -96 440795 -62 440811
rect -96 439803 -62 439819
rect 62 440795 96 440811
rect 62 439803 96 439819
rect -50 439735 -34 439769
rect 34 439735 50 439769
rect -50 439627 -34 439661
rect 34 439627 50 439661
rect -96 439577 -62 439593
rect -96 438585 -62 438601
rect 62 439577 96 439593
rect 62 438585 96 438601
rect -50 438517 -34 438551
rect 34 438517 50 438551
rect -50 438409 -34 438443
rect 34 438409 50 438443
rect -96 438359 -62 438375
rect -96 437367 -62 437383
rect 62 438359 96 438375
rect 62 437367 96 437383
rect -50 437299 -34 437333
rect 34 437299 50 437333
rect -50 437191 -34 437225
rect 34 437191 50 437225
rect -96 437141 -62 437157
rect -96 436149 -62 436165
rect 62 437141 96 437157
rect 62 436149 96 436165
rect -50 436081 -34 436115
rect 34 436081 50 436115
rect -50 435973 -34 436007
rect 34 435973 50 436007
rect -96 435923 -62 435939
rect -96 434931 -62 434947
rect 62 435923 96 435939
rect 62 434931 96 434947
rect -50 434863 -34 434897
rect 34 434863 50 434897
rect -50 434755 -34 434789
rect 34 434755 50 434789
rect -96 434705 -62 434721
rect -96 433713 -62 433729
rect 62 434705 96 434721
rect 62 433713 96 433729
rect -50 433645 -34 433679
rect 34 433645 50 433679
rect -50 433537 -34 433571
rect 34 433537 50 433571
rect -96 433487 -62 433503
rect -96 432495 -62 432511
rect 62 433487 96 433503
rect 62 432495 96 432511
rect -50 432427 -34 432461
rect 34 432427 50 432461
rect -50 432319 -34 432353
rect 34 432319 50 432353
rect -96 432269 -62 432285
rect -96 431277 -62 431293
rect 62 432269 96 432285
rect 62 431277 96 431293
rect -50 431209 -34 431243
rect 34 431209 50 431243
rect -50 431101 -34 431135
rect 34 431101 50 431135
rect -96 431051 -62 431067
rect -96 430059 -62 430075
rect 62 431051 96 431067
rect 62 430059 96 430075
rect -50 429991 -34 430025
rect 34 429991 50 430025
rect -50 429883 -34 429917
rect 34 429883 50 429917
rect -96 429833 -62 429849
rect -96 428841 -62 428857
rect 62 429833 96 429849
rect 62 428841 96 428857
rect -50 428773 -34 428807
rect 34 428773 50 428807
rect -50 428665 -34 428699
rect 34 428665 50 428699
rect -96 428615 -62 428631
rect -96 427623 -62 427639
rect 62 428615 96 428631
rect 62 427623 96 427639
rect -50 427555 -34 427589
rect 34 427555 50 427589
rect -50 427447 -34 427481
rect 34 427447 50 427481
rect -96 427397 -62 427413
rect -96 426405 -62 426421
rect 62 427397 96 427413
rect 62 426405 96 426421
rect -50 426337 -34 426371
rect 34 426337 50 426371
rect -50 426229 -34 426263
rect 34 426229 50 426263
rect -96 426179 -62 426195
rect -96 425187 -62 425203
rect 62 426179 96 426195
rect 62 425187 96 425203
rect -50 425119 -34 425153
rect 34 425119 50 425153
rect -50 425011 -34 425045
rect 34 425011 50 425045
rect -96 424961 -62 424977
rect -96 423969 -62 423985
rect 62 424961 96 424977
rect 62 423969 96 423985
rect -50 423901 -34 423935
rect 34 423901 50 423935
rect -50 423793 -34 423827
rect 34 423793 50 423827
rect -96 423743 -62 423759
rect -96 422751 -62 422767
rect 62 423743 96 423759
rect 62 422751 96 422767
rect -50 422683 -34 422717
rect 34 422683 50 422717
rect -50 422575 -34 422609
rect 34 422575 50 422609
rect -96 422525 -62 422541
rect -96 421533 -62 421549
rect 62 422525 96 422541
rect 62 421533 96 421549
rect -50 421465 -34 421499
rect 34 421465 50 421499
rect -50 421357 -34 421391
rect 34 421357 50 421391
rect -96 421307 -62 421323
rect -96 420315 -62 420331
rect 62 421307 96 421323
rect 62 420315 96 420331
rect -50 420247 -34 420281
rect 34 420247 50 420281
rect -50 420139 -34 420173
rect 34 420139 50 420173
rect -96 420089 -62 420105
rect -96 419097 -62 419113
rect 62 420089 96 420105
rect 62 419097 96 419113
rect -50 419029 -34 419063
rect 34 419029 50 419063
rect -50 418921 -34 418955
rect 34 418921 50 418955
rect -96 418871 -62 418887
rect -96 417879 -62 417895
rect 62 418871 96 418887
rect 62 417879 96 417895
rect -50 417811 -34 417845
rect 34 417811 50 417845
rect -50 417703 -34 417737
rect 34 417703 50 417737
rect -96 417653 -62 417669
rect -96 416661 -62 416677
rect 62 417653 96 417669
rect 62 416661 96 416677
rect -50 416593 -34 416627
rect 34 416593 50 416627
rect -50 416485 -34 416519
rect 34 416485 50 416519
rect -96 416435 -62 416451
rect -96 415443 -62 415459
rect 62 416435 96 416451
rect 62 415443 96 415459
rect -50 415375 -34 415409
rect 34 415375 50 415409
rect -50 415267 -34 415301
rect 34 415267 50 415301
rect -96 415217 -62 415233
rect -96 414225 -62 414241
rect 62 415217 96 415233
rect 62 414225 96 414241
rect -50 414157 -34 414191
rect 34 414157 50 414191
rect -50 414049 -34 414083
rect 34 414049 50 414083
rect -96 413999 -62 414015
rect -96 413007 -62 413023
rect 62 413999 96 414015
rect 62 413007 96 413023
rect -50 412939 -34 412973
rect 34 412939 50 412973
rect -50 412831 -34 412865
rect 34 412831 50 412865
rect -96 412781 -62 412797
rect -96 411789 -62 411805
rect 62 412781 96 412797
rect 62 411789 96 411805
rect -50 411721 -34 411755
rect 34 411721 50 411755
rect -50 411613 -34 411647
rect 34 411613 50 411647
rect -96 411563 -62 411579
rect -96 410571 -62 410587
rect 62 411563 96 411579
rect 62 410571 96 410587
rect -50 410503 -34 410537
rect 34 410503 50 410537
rect -50 410395 -34 410429
rect 34 410395 50 410429
rect -96 410345 -62 410361
rect -96 409353 -62 409369
rect 62 410345 96 410361
rect 62 409353 96 409369
rect -50 409285 -34 409319
rect 34 409285 50 409319
rect -50 409177 -34 409211
rect 34 409177 50 409211
rect -96 409127 -62 409143
rect -96 408135 -62 408151
rect 62 409127 96 409143
rect 62 408135 96 408151
rect -50 408067 -34 408101
rect 34 408067 50 408101
rect -50 407959 -34 407993
rect 34 407959 50 407993
rect -96 407909 -62 407925
rect -96 406917 -62 406933
rect 62 407909 96 407925
rect 62 406917 96 406933
rect -50 406849 -34 406883
rect 34 406849 50 406883
rect -50 406741 -34 406775
rect 34 406741 50 406775
rect -96 406691 -62 406707
rect -96 405699 -62 405715
rect 62 406691 96 406707
rect 62 405699 96 405715
rect -50 405631 -34 405665
rect 34 405631 50 405665
rect -50 405523 -34 405557
rect 34 405523 50 405557
rect -96 405473 -62 405489
rect -96 404481 -62 404497
rect 62 405473 96 405489
rect 62 404481 96 404497
rect -50 404413 -34 404447
rect 34 404413 50 404447
rect -50 404305 -34 404339
rect 34 404305 50 404339
rect -96 404255 -62 404271
rect -96 403263 -62 403279
rect 62 404255 96 404271
rect 62 403263 96 403279
rect -50 403195 -34 403229
rect 34 403195 50 403229
rect -50 403087 -34 403121
rect 34 403087 50 403121
rect -96 403037 -62 403053
rect -96 402045 -62 402061
rect 62 403037 96 403053
rect 62 402045 96 402061
rect -50 401977 -34 402011
rect 34 401977 50 402011
rect -50 401869 -34 401903
rect 34 401869 50 401903
rect -96 401819 -62 401835
rect -96 400827 -62 400843
rect 62 401819 96 401835
rect 62 400827 96 400843
rect -50 400759 -34 400793
rect 34 400759 50 400793
rect -50 400651 -34 400685
rect 34 400651 50 400685
rect -96 400601 -62 400617
rect -96 399609 -62 399625
rect 62 400601 96 400617
rect 62 399609 96 399625
rect -50 399541 -34 399575
rect 34 399541 50 399575
rect -50 399433 -34 399467
rect 34 399433 50 399467
rect -96 399383 -62 399399
rect -96 398391 -62 398407
rect 62 399383 96 399399
rect 62 398391 96 398407
rect -50 398323 -34 398357
rect 34 398323 50 398357
rect -50 398215 -34 398249
rect 34 398215 50 398249
rect -96 398165 -62 398181
rect -96 397173 -62 397189
rect 62 398165 96 398181
rect 62 397173 96 397189
rect -50 397105 -34 397139
rect 34 397105 50 397139
rect -50 396997 -34 397031
rect 34 396997 50 397031
rect -96 396947 -62 396963
rect -96 395955 -62 395971
rect 62 396947 96 396963
rect 62 395955 96 395971
rect -50 395887 -34 395921
rect 34 395887 50 395921
rect -50 395779 -34 395813
rect 34 395779 50 395813
rect -96 395729 -62 395745
rect -96 394737 -62 394753
rect 62 395729 96 395745
rect 62 394737 96 394753
rect -50 394669 -34 394703
rect 34 394669 50 394703
rect -50 394561 -34 394595
rect 34 394561 50 394595
rect -96 394511 -62 394527
rect -96 393519 -62 393535
rect 62 394511 96 394527
rect 62 393519 96 393535
rect -50 393451 -34 393485
rect 34 393451 50 393485
rect -50 393343 -34 393377
rect 34 393343 50 393377
rect -96 393293 -62 393309
rect -96 392301 -62 392317
rect 62 393293 96 393309
rect 62 392301 96 392317
rect -50 392233 -34 392267
rect 34 392233 50 392267
rect -50 392125 -34 392159
rect 34 392125 50 392159
rect -96 392075 -62 392091
rect -96 391083 -62 391099
rect 62 392075 96 392091
rect 62 391083 96 391099
rect -50 391015 -34 391049
rect 34 391015 50 391049
rect -50 390907 -34 390941
rect 34 390907 50 390941
rect -96 390857 -62 390873
rect -96 389865 -62 389881
rect 62 390857 96 390873
rect 62 389865 96 389881
rect -50 389797 -34 389831
rect 34 389797 50 389831
rect -50 389689 -34 389723
rect 34 389689 50 389723
rect -96 389639 -62 389655
rect -96 388647 -62 388663
rect 62 389639 96 389655
rect 62 388647 96 388663
rect -50 388579 -34 388613
rect 34 388579 50 388613
rect -50 388471 -34 388505
rect 34 388471 50 388505
rect -96 388421 -62 388437
rect -96 387429 -62 387445
rect 62 388421 96 388437
rect 62 387429 96 387445
rect -50 387361 -34 387395
rect 34 387361 50 387395
rect -50 387253 -34 387287
rect 34 387253 50 387287
rect -96 387203 -62 387219
rect -96 386211 -62 386227
rect 62 387203 96 387219
rect 62 386211 96 386227
rect -50 386143 -34 386177
rect 34 386143 50 386177
rect -50 386035 -34 386069
rect 34 386035 50 386069
rect -96 385985 -62 386001
rect -96 384993 -62 385009
rect 62 385985 96 386001
rect 62 384993 96 385009
rect -50 384925 -34 384959
rect 34 384925 50 384959
rect -50 384817 -34 384851
rect 34 384817 50 384851
rect -96 384767 -62 384783
rect -96 383775 -62 383791
rect 62 384767 96 384783
rect 62 383775 96 383791
rect -50 383707 -34 383741
rect 34 383707 50 383741
rect -50 383599 -34 383633
rect 34 383599 50 383633
rect -96 383549 -62 383565
rect -96 382557 -62 382573
rect 62 383549 96 383565
rect 62 382557 96 382573
rect -50 382489 -34 382523
rect 34 382489 50 382523
rect -50 382381 -34 382415
rect 34 382381 50 382415
rect -96 382331 -62 382347
rect -96 381339 -62 381355
rect 62 382331 96 382347
rect 62 381339 96 381355
rect -50 381271 -34 381305
rect 34 381271 50 381305
rect -50 381163 -34 381197
rect 34 381163 50 381197
rect -96 381113 -62 381129
rect -96 380121 -62 380137
rect 62 381113 96 381129
rect 62 380121 96 380137
rect -50 380053 -34 380087
rect 34 380053 50 380087
rect -50 379945 -34 379979
rect 34 379945 50 379979
rect -96 379895 -62 379911
rect -96 378903 -62 378919
rect 62 379895 96 379911
rect 62 378903 96 378919
rect -50 378835 -34 378869
rect 34 378835 50 378869
rect -50 378727 -34 378761
rect 34 378727 50 378761
rect -96 378677 -62 378693
rect -96 377685 -62 377701
rect 62 378677 96 378693
rect 62 377685 96 377701
rect -50 377617 -34 377651
rect 34 377617 50 377651
rect -50 377509 -34 377543
rect 34 377509 50 377543
rect -96 377459 -62 377475
rect -96 376467 -62 376483
rect 62 377459 96 377475
rect 62 376467 96 376483
rect -50 376399 -34 376433
rect 34 376399 50 376433
rect -50 376291 -34 376325
rect 34 376291 50 376325
rect -96 376241 -62 376257
rect -96 375249 -62 375265
rect 62 376241 96 376257
rect 62 375249 96 375265
rect -50 375181 -34 375215
rect 34 375181 50 375215
rect -50 375073 -34 375107
rect 34 375073 50 375107
rect -96 375023 -62 375039
rect -96 374031 -62 374047
rect 62 375023 96 375039
rect 62 374031 96 374047
rect -50 373963 -34 373997
rect 34 373963 50 373997
rect -50 373855 -34 373889
rect 34 373855 50 373889
rect -96 373805 -62 373821
rect -96 372813 -62 372829
rect 62 373805 96 373821
rect 62 372813 96 372829
rect -50 372745 -34 372779
rect 34 372745 50 372779
rect -50 372637 -34 372671
rect 34 372637 50 372671
rect -96 372587 -62 372603
rect -96 371595 -62 371611
rect 62 372587 96 372603
rect 62 371595 96 371611
rect -50 371527 -34 371561
rect 34 371527 50 371561
rect -50 371419 -34 371453
rect 34 371419 50 371453
rect -96 371369 -62 371385
rect -96 370377 -62 370393
rect 62 371369 96 371385
rect 62 370377 96 370393
rect -50 370309 -34 370343
rect 34 370309 50 370343
rect -50 370201 -34 370235
rect 34 370201 50 370235
rect -96 370151 -62 370167
rect -96 369159 -62 369175
rect 62 370151 96 370167
rect 62 369159 96 369175
rect -50 369091 -34 369125
rect 34 369091 50 369125
rect -50 368983 -34 369017
rect 34 368983 50 369017
rect -96 368933 -62 368949
rect -96 367941 -62 367957
rect 62 368933 96 368949
rect 62 367941 96 367957
rect -50 367873 -34 367907
rect 34 367873 50 367907
rect -50 367765 -34 367799
rect 34 367765 50 367799
rect -96 367715 -62 367731
rect -96 366723 -62 366739
rect 62 367715 96 367731
rect 62 366723 96 366739
rect -50 366655 -34 366689
rect 34 366655 50 366689
rect -50 366547 -34 366581
rect 34 366547 50 366581
rect -96 366497 -62 366513
rect -96 365505 -62 365521
rect 62 366497 96 366513
rect 62 365505 96 365521
rect -50 365437 -34 365471
rect 34 365437 50 365471
rect -50 365329 -34 365363
rect 34 365329 50 365363
rect -96 365279 -62 365295
rect -96 364287 -62 364303
rect 62 365279 96 365295
rect 62 364287 96 364303
rect -50 364219 -34 364253
rect 34 364219 50 364253
rect -50 364111 -34 364145
rect 34 364111 50 364145
rect -96 364061 -62 364077
rect -96 363069 -62 363085
rect 62 364061 96 364077
rect 62 363069 96 363085
rect -50 363001 -34 363035
rect 34 363001 50 363035
rect -50 362893 -34 362927
rect 34 362893 50 362927
rect -96 362843 -62 362859
rect -96 361851 -62 361867
rect 62 362843 96 362859
rect 62 361851 96 361867
rect -50 361783 -34 361817
rect 34 361783 50 361817
rect -50 361675 -34 361709
rect 34 361675 50 361709
rect -96 361625 -62 361641
rect -96 360633 -62 360649
rect 62 361625 96 361641
rect 62 360633 96 360649
rect -50 360565 -34 360599
rect 34 360565 50 360599
rect -50 360457 -34 360491
rect 34 360457 50 360491
rect -96 360407 -62 360423
rect -96 359415 -62 359431
rect 62 360407 96 360423
rect 62 359415 96 359431
rect -50 359347 -34 359381
rect 34 359347 50 359381
rect -50 359239 -34 359273
rect 34 359239 50 359273
rect -96 359189 -62 359205
rect -96 358197 -62 358213
rect 62 359189 96 359205
rect 62 358197 96 358213
rect -50 358129 -34 358163
rect 34 358129 50 358163
rect -50 358021 -34 358055
rect 34 358021 50 358055
rect -96 357971 -62 357987
rect -96 356979 -62 356995
rect 62 357971 96 357987
rect 62 356979 96 356995
rect -50 356911 -34 356945
rect 34 356911 50 356945
rect -50 356803 -34 356837
rect 34 356803 50 356837
rect -96 356753 -62 356769
rect -96 355761 -62 355777
rect 62 356753 96 356769
rect 62 355761 96 355777
rect -50 355693 -34 355727
rect 34 355693 50 355727
rect -50 355585 -34 355619
rect 34 355585 50 355619
rect -96 355535 -62 355551
rect -96 354543 -62 354559
rect 62 355535 96 355551
rect 62 354543 96 354559
rect -50 354475 -34 354509
rect 34 354475 50 354509
rect -50 354367 -34 354401
rect 34 354367 50 354401
rect -96 354317 -62 354333
rect -96 353325 -62 353341
rect 62 354317 96 354333
rect 62 353325 96 353341
rect -50 353257 -34 353291
rect 34 353257 50 353291
rect -50 353149 -34 353183
rect 34 353149 50 353183
rect -96 353099 -62 353115
rect -96 352107 -62 352123
rect 62 353099 96 353115
rect 62 352107 96 352123
rect -50 352039 -34 352073
rect 34 352039 50 352073
rect -50 351931 -34 351965
rect 34 351931 50 351965
rect -96 351881 -62 351897
rect -96 350889 -62 350905
rect 62 351881 96 351897
rect 62 350889 96 350905
rect -50 350821 -34 350855
rect 34 350821 50 350855
rect -50 350713 -34 350747
rect 34 350713 50 350747
rect -96 350663 -62 350679
rect -96 349671 -62 349687
rect 62 350663 96 350679
rect 62 349671 96 349687
rect -50 349603 -34 349637
rect 34 349603 50 349637
rect -50 349495 -34 349529
rect 34 349495 50 349529
rect -96 349445 -62 349461
rect -96 348453 -62 348469
rect 62 349445 96 349461
rect 62 348453 96 348469
rect -50 348385 -34 348419
rect 34 348385 50 348419
rect -50 348277 -34 348311
rect 34 348277 50 348311
rect -96 348227 -62 348243
rect -96 347235 -62 347251
rect 62 348227 96 348243
rect 62 347235 96 347251
rect -50 347167 -34 347201
rect 34 347167 50 347201
rect -50 347059 -34 347093
rect 34 347059 50 347093
rect -96 347009 -62 347025
rect -96 346017 -62 346033
rect 62 347009 96 347025
rect 62 346017 96 346033
rect -50 345949 -34 345983
rect 34 345949 50 345983
rect -50 345841 -34 345875
rect 34 345841 50 345875
rect -96 345791 -62 345807
rect -96 344799 -62 344815
rect 62 345791 96 345807
rect 62 344799 96 344815
rect -50 344731 -34 344765
rect 34 344731 50 344765
rect -50 344623 -34 344657
rect 34 344623 50 344657
rect -96 344573 -62 344589
rect -96 343581 -62 343597
rect 62 344573 96 344589
rect 62 343581 96 343597
rect -50 343513 -34 343547
rect 34 343513 50 343547
rect -50 343405 -34 343439
rect 34 343405 50 343439
rect -96 343355 -62 343371
rect -96 342363 -62 342379
rect 62 343355 96 343371
rect 62 342363 96 342379
rect -50 342295 -34 342329
rect 34 342295 50 342329
rect -50 342187 -34 342221
rect 34 342187 50 342221
rect -96 342137 -62 342153
rect -96 341145 -62 341161
rect 62 342137 96 342153
rect 62 341145 96 341161
rect -50 341077 -34 341111
rect 34 341077 50 341111
rect -50 340969 -34 341003
rect 34 340969 50 341003
rect -96 340919 -62 340935
rect -96 339927 -62 339943
rect 62 340919 96 340935
rect 62 339927 96 339943
rect -50 339859 -34 339893
rect 34 339859 50 339893
rect -50 339751 -34 339785
rect 34 339751 50 339785
rect -96 339701 -62 339717
rect -96 338709 -62 338725
rect 62 339701 96 339717
rect 62 338709 96 338725
rect -50 338641 -34 338675
rect 34 338641 50 338675
rect -50 338533 -34 338567
rect 34 338533 50 338567
rect -96 338483 -62 338499
rect -96 337491 -62 337507
rect 62 338483 96 338499
rect 62 337491 96 337507
rect -50 337423 -34 337457
rect 34 337423 50 337457
rect -50 337315 -34 337349
rect 34 337315 50 337349
rect -96 337265 -62 337281
rect -96 336273 -62 336289
rect 62 337265 96 337281
rect 62 336273 96 336289
rect -50 336205 -34 336239
rect 34 336205 50 336239
rect -50 336097 -34 336131
rect 34 336097 50 336131
rect -96 336047 -62 336063
rect -96 335055 -62 335071
rect 62 336047 96 336063
rect 62 335055 96 335071
rect -50 334987 -34 335021
rect 34 334987 50 335021
rect -50 334879 -34 334913
rect 34 334879 50 334913
rect -96 334829 -62 334845
rect -96 333837 -62 333853
rect 62 334829 96 334845
rect 62 333837 96 333853
rect -50 333769 -34 333803
rect 34 333769 50 333803
rect -50 333661 -34 333695
rect 34 333661 50 333695
rect -96 333611 -62 333627
rect -96 332619 -62 332635
rect 62 333611 96 333627
rect 62 332619 96 332635
rect -50 332551 -34 332585
rect 34 332551 50 332585
rect -50 332443 -34 332477
rect 34 332443 50 332477
rect -96 332393 -62 332409
rect -96 331401 -62 331417
rect 62 332393 96 332409
rect 62 331401 96 331417
rect -50 331333 -34 331367
rect 34 331333 50 331367
rect -50 331225 -34 331259
rect 34 331225 50 331259
rect -96 331175 -62 331191
rect -96 330183 -62 330199
rect 62 331175 96 331191
rect 62 330183 96 330199
rect -50 330115 -34 330149
rect 34 330115 50 330149
rect -50 330007 -34 330041
rect 34 330007 50 330041
rect -96 329957 -62 329973
rect -96 328965 -62 328981
rect 62 329957 96 329973
rect 62 328965 96 328981
rect -50 328897 -34 328931
rect 34 328897 50 328931
rect -50 328789 -34 328823
rect 34 328789 50 328823
rect -96 328739 -62 328755
rect -96 327747 -62 327763
rect 62 328739 96 328755
rect 62 327747 96 327763
rect -50 327679 -34 327713
rect 34 327679 50 327713
rect -50 327571 -34 327605
rect 34 327571 50 327605
rect -96 327521 -62 327537
rect -96 326529 -62 326545
rect 62 327521 96 327537
rect 62 326529 96 326545
rect -50 326461 -34 326495
rect 34 326461 50 326495
rect -50 326353 -34 326387
rect 34 326353 50 326387
rect -96 326303 -62 326319
rect -96 325311 -62 325327
rect 62 326303 96 326319
rect 62 325311 96 325327
rect -50 325243 -34 325277
rect 34 325243 50 325277
rect -50 325135 -34 325169
rect 34 325135 50 325169
rect -96 325085 -62 325101
rect -96 324093 -62 324109
rect 62 325085 96 325101
rect 62 324093 96 324109
rect -50 324025 -34 324059
rect 34 324025 50 324059
rect -50 323917 -34 323951
rect 34 323917 50 323951
rect -96 323867 -62 323883
rect -96 322875 -62 322891
rect 62 323867 96 323883
rect 62 322875 96 322891
rect -50 322807 -34 322841
rect 34 322807 50 322841
rect -50 322699 -34 322733
rect 34 322699 50 322733
rect -96 322649 -62 322665
rect -96 321657 -62 321673
rect 62 322649 96 322665
rect 62 321657 96 321673
rect -50 321589 -34 321623
rect 34 321589 50 321623
rect -50 321481 -34 321515
rect 34 321481 50 321515
rect -96 321431 -62 321447
rect -96 320439 -62 320455
rect 62 321431 96 321447
rect 62 320439 96 320455
rect -50 320371 -34 320405
rect 34 320371 50 320405
rect -50 320263 -34 320297
rect 34 320263 50 320297
rect -96 320213 -62 320229
rect -96 319221 -62 319237
rect 62 320213 96 320229
rect 62 319221 96 319237
rect -50 319153 -34 319187
rect 34 319153 50 319187
rect -50 319045 -34 319079
rect 34 319045 50 319079
rect -96 318995 -62 319011
rect -96 318003 -62 318019
rect 62 318995 96 319011
rect 62 318003 96 318019
rect -50 317935 -34 317969
rect 34 317935 50 317969
rect -50 317827 -34 317861
rect 34 317827 50 317861
rect -96 317777 -62 317793
rect -96 316785 -62 316801
rect 62 317777 96 317793
rect 62 316785 96 316801
rect -50 316717 -34 316751
rect 34 316717 50 316751
rect -50 316609 -34 316643
rect 34 316609 50 316643
rect -96 316559 -62 316575
rect -96 315567 -62 315583
rect 62 316559 96 316575
rect 62 315567 96 315583
rect -50 315499 -34 315533
rect 34 315499 50 315533
rect -50 315391 -34 315425
rect 34 315391 50 315425
rect -96 315341 -62 315357
rect -96 314349 -62 314365
rect 62 315341 96 315357
rect 62 314349 96 314365
rect -50 314281 -34 314315
rect 34 314281 50 314315
rect -50 314173 -34 314207
rect 34 314173 50 314207
rect -96 314123 -62 314139
rect -96 313131 -62 313147
rect 62 314123 96 314139
rect 62 313131 96 313147
rect -50 313063 -34 313097
rect 34 313063 50 313097
rect -50 312955 -34 312989
rect 34 312955 50 312989
rect -96 312905 -62 312921
rect -96 311913 -62 311929
rect 62 312905 96 312921
rect 62 311913 96 311929
rect -50 311845 -34 311879
rect 34 311845 50 311879
rect -50 311737 -34 311771
rect 34 311737 50 311771
rect -96 311687 -62 311703
rect -96 310695 -62 310711
rect 62 311687 96 311703
rect 62 310695 96 310711
rect -50 310627 -34 310661
rect 34 310627 50 310661
rect -50 310519 -34 310553
rect 34 310519 50 310553
rect -96 310469 -62 310485
rect -96 309477 -62 309493
rect 62 310469 96 310485
rect 62 309477 96 309493
rect -50 309409 -34 309443
rect 34 309409 50 309443
rect -50 309301 -34 309335
rect 34 309301 50 309335
rect -96 309251 -62 309267
rect -96 308259 -62 308275
rect 62 309251 96 309267
rect 62 308259 96 308275
rect -50 308191 -34 308225
rect 34 308191 50 308225
rect -50 308083 -34 308117
rect 34 308083 50 308117
rect -96 308033 -62 308049
rect -96 307041 -62 307057
rect 62 308033 96 308049
rect 62 307041 96 307057
rect -50 306973 -34 307007
rect 34 306973 50 307007
rect -50 306865 -34 306899
rect 34 306865 50 306899
rect -96 306815 -62 306831
rect -96 305823 -62 305839
rect 62 306815 96 306831
rect 62 305823 96 305839
rect -50 305755 -34 305789
rect 34 305755 50 305789
rect -50 305647 -34 305681
rect 34 305647 50 305681
rect -96 305597 -62 305613
rect -96 304605 -62 304621
rect 62 305597 96 305613
rect 62 304605 96 304621
rect -50 304537 -34 304571
rect 34 304537 50 304571
rect -50 304429 -34 304463
rect 34 304429 50 304463
rect -96 304379 -62 304395
rect -96 303387 -62 303403
rect 62 304379 96 304395
rect 62 303387 96 303403
rect -50 303319 -34 303353
rect 34 303319 50 303353
rect -50 303211 -34 303245
rect 34 303211 50 303245
rect -96 303161 -62 303177
rect -96 302169 -62 302185
rect 62 303161 96 303177
rect 62 302169 96 302185
rect -50 302101 -34 302135
rect 34 302101 50 302135
rect -50 301993 -34 302027
rect 34 301993 50 302027
rect -96 301943 -62 301959
rect -96 300951 -62 300967
rect 62 301943 96 301959
rect 62 300951 96 300967
rect -50 300883 -34 300917
rect 34 300883 50 300917
rect -50 300775 -34 300809
rect 34 300775 50 300809
rect -96 300725 -62 300741
rect -96 299733 -62 299749
rect 62 300725 96 300741
rect 62 299733 96 299749
rect -50 299665 -34 299699
rect 34 299665 50 299699
rect -50 299557 -34 299591
rect 34 299557 50 299591
rect -96 299507 -62 299523
rect -96 298515 -62 298531
rect 62 299507 96 299523
rect 62 298515 96 298531
rect -50 298447 -34 298481
rect 34 298447 50 298481
rect -50 298339 -34 298373
rect 34 298339 50 298373
rect -96 298289 -62 298305
rect -96 297297 -62 297313
rect 62 298289 96 298305
rect 62 297297 96 297313
rect -50 297229 -34 297263
rect 34 297229 50 297263
rect -50 297121 -34 297155
rect 34 297121 50 297155
rect -96 297071 -62 297087
rect -96 296079 -62 296095
rect 62 297071 96 297087
rect 62 296079 96 296095
rect -50 296011 -34 296045
rect 34 296011 50 296045
rect -50 295903 -34 295937
rect 34 295903 50 295937
rect -96 295853 -62 295869
rect -96 294861 -62 294877
rect 62 295853 96 295869
rect 62 294861 96 294877
rect -50 294793 -34 294827
rect 34 294793 50 294827
rect -50 294685 -34 294719
rect 34 294685 50 294719
rect -96 294635 -62 294651
rect -96 293643 -62 293659
rect 62 294635 96 294651
rect 62 293643 96 293659
rect -50 293575 -34 293609
rect 34 293575 50 293609
rect -50 293467 -34 293501
rect 34 293467 50 293501
rect -96 293417 -62 293433
rect -96 292425 -62 292441
rect 62 293417 96 293433
rect 62 292425 96 292441
rect -50 292357 -34 292391
rect 34 292357 50 292391
rect -50 292249 -34 292283
rect 34 292249 50 292283
rect -96 292199 -62 292215
rect -96 291207 -62 291223
rect 62 292199 96 292215
rect 62 291207 96 291223
rect -50 291139 -34 291173
rect 34 291139 50 291173
rect -50 291031 -34 291065
rect 34 291031 50 291065
rect -96 290981 -62 290997
rect -96 289989 -62 290005
rect 62 290981 96 290997
rect 62 289989 96 290005
rect -50 289921 -34 289955
rect 34 289921 50 289955
rect -50 289813 -34 289847
rect 34 289813 50 289847
rect -96 289763 -62 289779
rect -96 288771 -62 288787
rect 62 289763 96 289779
rect 62 288771 96 288787
rect -50 288703 -34 288737
rect 34 288703 50 288737
rect -50 288595 -34 288629
rect 34 288595 50 288629
rect -96 288545 -62 288561
rect -96 287553 -62 287569
rect 62 288545 96 288561
rect 62 287553 96 287569
rect -50 287485 -34 287519
rect 34 287485 50 287519
rect -50 287377 -34 287411
rect 34 287377 50 287411
rect -96 287327 -62 287343
rect -96 286335 -62 286351
rect 62 287327 96 287343
rect 62 286335 96 286351
rect -50 286267 -34 286301
rect 34 286267 50 286301
rect -50 286159 -34 286193
rect 34 286159 50 286193
rect -96 286109 -62 286125
rect -96 285117 -62 285133
rect 62 286109 96 286125
rect 62 285117 96 285133
rect -50 285049 -34 285083
rect 34 285049 50 285083
rect -50 284941 -34 284975
rect 34 284941 50 284975
rect -96 284891 -62 284907
rect -96 283899 -62 283915
rect 62 284891 96 284907
rect 62 283899 96 283915
rect -50 283831 -34 283865
rect 34 283831 50 283865
rect -50 283723 -34 283757
rect 34 283723 50 283757
rect -96 283673 -62 283689
rect -96 282681 -62 282697
rect 62 283673 96 283689
rect 62 282681 96 282697
rect -50 282613 -34 282647
rect 34 282613 50 282647
rect -50 282505 -34 282539
rect 34 282505 50 282539
rect -96 282455 -62 282471
rect -96 281463 -62 281479
rect 62 282455 96 282471
rect 62 281463 96 281479
rect -50 281395 -34 281429
rect 34 281395 50 281429
rect -50 281287 -34 281321
rect 34 281287 50 281321
rect -96 281237 -62 281253
rect -96 280245 -62 280261
rect 62 281237 96 281253
rect 62 280245 96 280261
rect -50 280177 -34 280211
rect 34 280177 50 280211
rect -50 280069 -34 280103
rect 34 280069 50 280103
rect -96 280019 -62 280035
rect -96 279027 -62 279043
rect 62 280019 96 280035
rect 62 279027 96 279043
rect -50 278959 -34 278993
rect 34 278959 50 278993
rect -50 278851 -34 278885
rect 34 278851 50 278885
rect -96 278801 -62 278817
rect -96 277809 -62 277825
rect 62 278801 96 278817
rect 62 277809 96 277825
rect -50 277741 -34 277775
rect 34 277741 50 277775
rect -50 277633 -34 277667
rect 34 277633 50 277667
rect -96 277583 -62 277599
rect -96 276591 -62 276607
rect 62 277583 96 277599
rect 62 276591 96 276607
rect -50 276523 -34 276557
rect 34 276523 50 276557
rect -50 276415 -34 276449
rect 34 276415 50 276449
rect -96 276365 -62 276381
rect -96 275373 -62 275389
rect 62 276365 96 276381
rect 62 275373 96 275389
rect -50 275305 -34 275339
rect 34 275305 50 275339
rect -50 275197 -34 275231
rect 34 275197 50 275231
rect -96 275147 -62 275163
rect -96 274155 -62 274171
rect 62 275147 96 275163
rect 62 274155 96 274171
rect -50 274087 -34 274121
rect 34 274087 50 274121
rect -50 273979 -34 274013
rect 34 273979 50 274013
rect -96 273929 -62 273945
rect -96 272937 -62 272953
rect 62 273929 96 273945
rect 62 272937 96 272953
rect -50 272869 -34 272903
rect 34 272869 50 272903
rect -50 272761 -34 272795
rect 34 272761 50 272795
rect -96 272711 -62 272727
rect -96 271719 -62 271735
rect 62 272711 96 272727
rect 62 271719 96 271735
rect -50 271651 -34 271685
rect 34 271651 50 271685
rect -50 271543 -34 271577
rect 34 271543 50 271577
rect -96 271493 -62 271509
rect -96 270501 -62 270517
rect 62 271493 96 271509
rect 62 270501 96 270517
rect -50 270433 -34 270467
rect 34 270433 50 270467
rect -50 270325 -34 270359
rect 34 270325 50 270359
rect -96 270275 -62 270291
rect -96 269283 -62 269299
rect 62 270275 96 270291
rect 62 269283 96 269299
rect -50 269215 -34 269249
rect 34 269215 50 269249
rect -50 269107 -34 269141
rect 34 269107 50 269141
rect -96 269057 -62 269073
rect -96 268065 -62 268081
rect 62 269057 96 269073
rect 62 268065 96 268081
rect -50 267997 -34 268031
rect 34 267997 50 268031
rect -50 267889 -34 267923
rect 34 267889 50 267923
rect -96 267839 -62 267855
rect -96 266847 -62 266863
rect 62 267839 96 267855
rect 62 266847 96 266863
rect -50 266779 -34 266813
rect 34 266779 50 266813
rect -50 266671 -34 266705
rect 34 266671 50 266705
rect -96 266621 -62 266637
rect -96 265629 -62 265645
rect 62 266621 96 266637
rect 62 265629 96 265645
rect -50 265561 -34 265595
rect 34 265561 50 265595
rect -50 265453 -34 265487
rect 34 265453 50 265487
rect -96 265403 -62 265419
rect -96 264411 -62 264427
rect 62 265403 96 265419
rect 62 264411 96 264427
rect -50 264343 -34 264377
rect 34 264343 50 264377
rect -50 264235 -34 264269
rect 34 264235 50 264269
rect -96 264185 -62 264201
rect -96 263193 -62 263209
rect 62 264185 96 264201
rect 62 263193 96 263209
rect -50 263125 -34 263159
rect 34 263125 50 263159
rect -50 263017 -34 263051
rect 34 263017 50 263051
rect -96 262967 -62 262983
rect -96 261975 -62 261991
rect 62 262967 96 262983
rect 62 261975 96 261991
rect -50 261907 -34 261941
rect 34 261907 50 261941
rect -50 261799 -34 261833
rect 34 261799 50 261833
rect -96 261749 -62 261765
rect -96 260757 -62 260773
rect 62 261749 96 261765
rect 62 260757 96 260773
rect -50 260689 -34 260723
rect 34 260689 50 260723
rect -50 260581 -34 260615
rect 34 260581 50 260615
rect -96 260531 -62 260547
rect -96 259539 -62 259555
rect 62 260531 96 260547
rect 62 259539 96 259555
rect -50 259471 -34 259505
rect 34 259471 50 259505
rect -50 259363 -34 259397
rect 34 259363 50 259397
rect -96 259313 -62 259329
rect -96 258321 -62 258337
rect 62 259313 96 259329
rect 62 258321 96 258337
rect -50 258253 -34 258287
rect 34 258253 50 258287
rect -50 258145 -34 258179
rect 34 258145 50 258179
rect -96 258095 -62 258111
rect -96 257103 -62 257119
rect 62 258095 96 258111
rect 62 257103 96 257119
rect -50 257035 -34 257069
rect 34 257035 50 257069
rect -50 256927 -34 256961
rect 34 256927 50 256961
rect -96 256877 -62 256893
rect -96 255885 -62 255901
rect 62 256877 96 256893
rect 62 255885 96 255901
rect -50 255817 -34 255851
rect 34 255817 50 255851
rect -50 255709 -34 255743
rect 34 255709 50 255743
rect -96 255659 -62 255675
rect -96 254667 -62 254683
rect 62 255659 96 255675
rect 62 254667 96 254683
rect -50 254599 -34 254633
rect 34 254599 50 254633
rect -50 254491 -34 254525
rect 34 254491 50 254525
rect -96 254441 -62 254457
rect -96 253449 -62 253465
rect 62 254441 96 254457
rect 62 253449 96 253465
rect -50 253381 -34 253415
rect 34 253381 50 253415
rect -50 253273 -34 253307
rect 34 253273 50 253307
rect -96 253223 -62 253239
rect -96 252231 -62 252247
rect 62 253223 96 253239
rect 62 252231 96 252247
rect -50 252163 -34 252197
rect 34 252163 50 252197
rect -50 252055 -34 252089
rect 34 252055 50 252089
rect -96 252005 -62 252021
rect -96 251013 -62 251029
rect 62 252005 96 252021
rect 62 251013 96 251029
rect -50 250945 -34 250979
rect 34 250945 50 250979
rect -50 250837 -34 250871
rect 34 250837 50 250871
rect -96 250787 -62 250803
rect -96 249795 -62 249811
rect 62 250787 96 250803
rect 62 249795 96 249811
rect -50 249727 -34 249761
rect 34 249727 50 249761
rect -50 249619 -34 249653
rect 34 249619 50 249653
rect -96 249569 -62 249585
rect -96 248577 -62 248593
rect 62 249569 96 249585
rect 62 248577 96 248593
rect -50 248509 -34 248543
rect 34 248509 50 248543
rect -50 248401 -34 248435
rect 34 248401 50 248435
rect -96 248351 -62 248367
rect -96 247359 -62 247375
rect 62 248351 96 248367
rect 62 247359 96 247375
rect -50 247291 -34 247325
rect 34 247291 50 247325
rect -50 247183 -34 247217
rect 34 247183 50 247217
rect -96 247133 -62 247149
rect -96 246141 -62 246157
rect 62 247133 96 247149
rect 62 246141 96 246157
rect -50 246073 -34 246107
rect 34 246073 50 246107
rect -50 245965 -34 245999
rect 34 245965 50 245999
rect -96 245915 -62 245931
rect -96 244923 -62 244939
rect 62 245915 96 245931
rect 62 244923 96 244939
rect -50 244855 -34 244889
rect 34 244855 50 244889
rect -50 244747 -34 244781
rect 34 244747 50 244781
rect -96 244697 -62 244713
rect -96 243705 -62 243721
rect 62 244697 96 244713
rect 62 243705 96 243721
rect -50 243637 -34 243671
rect 34 243637 50 243671
rect -50 243529 -34 243563
rect 34 243529 50 243563
rect -96 243479 -62 243495
rect -96 242487 -62 242503
rect 62 243479 96 243495
rect 62 242487 96 242503
rect -50 242419 -34 242453
rect 34 242419 50 242453
rect -50 242311 -34 242345
rect 34 242311 50 242345
rect -96 242261 -62 242277
rect -96 241269 -62 241285
rect 62 242261 96 242277
rect 62 241269 96 241285
rect -50 241201 -34 241235
rect 34 241201 50 241235
rect -50 241093 -34 241127
rect 34 241093 50 241127
rect -96 241043 -62 241059
rect -96 240051 -62 240067
rect 62 241043 96 241059
rect 62 240051 96 240067
rect -50 239983 -34 240017
rect 34 239983 50 240017
rect -50 239875 -34 239909
rect 34 239875 50 239909
rect -96 239825 -62 239841
rect -96 238833 -62 238849
rect 62 239825 96 239841
rect 62 238833 96 238849
rect -50 238765 -34 238799
rect 34 238765 50 238799
rect -50 238657 -34 238691
rect 34 238657 50 238691
rect -96 238607 -62 238623
rect -96 237615 -62 237631
rect 62 238607 96 238623
rect 62 237615 96 237631
rect -50 237547 -34 237581
rect 34 237547 50 237581
rect -50 237439 -34 237473
rect 34 237439 50 237473
rect -96 237389 -62 237405
rect -96 236397 -62 236413
rect 62 237389 96 237405
rect 62 236397 96 236413
rect -50 236329 -34 236363
rect 34 236329 50 236363
rect -50 236221 -34 236255
rect 34 236221 50 236255
rect -96 236171 -62 236187
rect -96 235179 -62 235195
rect 62 236171 96 236187
rect 62 235179 96 235195
rect -50 235111 -34 235145
rect 34 235111 50 235145
rect -50 235003 -34 235037
rect 34 235003 50 235037
rect -96 234953 -62 234969
rect -96 233961 -62 233977
rect 62 234953 96 234969
rect 62 233961 96 233977
rect -50 233893 -34 233927
rect 34 233893 50 233927
rect -50 233785 -34 233819
rect 34 233785 50 233819
rect -96 233735 -62 233751
rect -96 232743 -62 232759
rect 62 233735 96 233751
rect 62 232743 96 232759
rect -50 232675 -34 232709
rect 34 232675 50 232709
rect -50 232567 -34 232601
rect 34 232567 50 232601
rect -96 232517 -62 232533
rect -96 231525 -62 231541
rect 62 232517 96 232533
rect 62 231525 96 231541
rect -50 231457 -34 231491
rect 34 231457 50 231491
rect -50 231349 -34 231383
rect 34 231349 50 231383
rect -96 231299 -62 231315
rect -96 230307 -62 230323
rect 62 231299 96 231315
rect 62 230307 96 230323
rect -50 230239 -34 230273
rect 34 230239 50 230273
rect -50 230131 -34 230165
rect 34 230131 50 230165
rect -96 230081 -62 230097
rect -96 229089 -62 229105
rect 62 230081 96 230097
rect 62 229089 96 229105
rect -50 229021 -34 229055
rect 34 229021 50 229055
rect -50 228913 -34 228947
rect 34 228913 50 228947
rect -96 228863 -62 228879
rect -96 227871 -62 227887
rect 62 228863 96 228879
rect 62 227871 96 227887
rect -50 227803 -34 227837
rect 34 227803 50 227837
rect -50 227695 -34 227729
rect 34 227695 50 227729
rect -96 227645 -62 227661
rect -96 226653 -62 226669
rect 62 227645 96 227661
rect 62 226653 96 226669
rect -50 226585 -34 226619
rect 34 226585 50 226619
rect -50 226477 -34 226511
rect 34 226477 50 226511
rect -96 226427 -62 226443
rect -96 225435 -62 225451
rect 62 226427 96 226443
rect 62 225435 96 225451
rect -50 225367 -34 225401
rect 34 225367 50 225401
rect -50 225259 -34 225293
rect 34 225259 50 225293
rect -96 225209 -62 225225
rect -96 224217 -62 224233
rect 62 225209 96 225225
rect 62 224217 96 224233
rect -50 224149 -34 224183
rect 34 224149 50 224183
rect -50 224041 -34 224075
rect 34 224041 50 224075
rect -96 223991 -62 224007
rect -96 222999 -62 223015
rect 62 223991 96 224007
rect 62 222999 96 223015
rect -50 222931 -34 222965
rect 34 222931 50 222965
rect -50 222823 -34 222857
rect 34 222823 50 222857
rect -96 222773 -62 222789
rect -96 221781 -62 221797
rect 62 222773 96 222789
rect 62 221781 96 221797
rect -50 221713 -34 221747
rect 34 221713 50 221747
rect -50 221605 -34 221639
rect 34 221605 50 221639
rect -96 221555 -62 221571
rect -96 220563 -62 220579
rect 62 221555 96 221571
rect 62 220563 96 220579
rect -50 220495 -34 220529
rect 34 220495 50 220529
rect -50 220387 -34 220421
rect 34 220387 50 220421
rect -96 220337 -62 220353
rect -96 219345 -62 219361
rect 62 220337 96 220353
rect 62 219345 96 219361
rect -50 219277 -34 219311
rect 34 219277 50 219311
rect -50 219169 -34 219203
rect 34 219169 50 219203
rect -96 219119 -62 219135
rect -96 218127 -62 218143
rect 62 219119 96 219135
rect 62 218127 96 218143
rect -50 218059 -34 218093
rect 34 218059 50 218093
rect -50 217951 -34 217985
rect 34 217951 50 217985
rect -96 217901 -62 217917
rect -96 216909 -62 216925
rect 62 217901 96 217917
rect 62 216909 96 216925
rect -50 216841 -34 216875
rect 34 216841 50 216875
rect -50 216733 -34 216767
rect 34 216733 50 216767
rect -96 216683 -62 216699
rect -96 215691 -62 215707
rect 62 216683 96 216699
rect 62 215691 96 215707
rect -50 215623 -34 215657
rect 34 215623 50 215657
rect -50 215515 -34 215549
rect 34 215515 50 215549
rect -96 215465 -62 215481
rect -96 214473 -62 214489
rect 62 215465 96 215481
rect 62 214473 96 214489
rect -50 214405 -34 214439
rect 34 214405 50 214439
rect -50 214297 -34 214331
rect 34 214297 50 214331
rect -96 214247 -62 214263
rect -96 213255 -62 213271
rect 62 214247 96 214263
rect 62 213255 96 213271
rect -50 213187 -34 213221
rect 34 213187 50 213221
rect -50 213079 -34 213113
rect 34 213079 50 213113
rect -96 213029 -62 213045
rect -96 212037 -62 212053
rect 62 213029 96 213045
rect 62 212037 96 212053
rect -50 211969 -34 212003
rect 34 211969 50 212003
rect -50 211861 -34 211895
rect 34 211861 50 211895
rect -96 211811 -62 211827
rect -96 210819 -62 210835
rect 62 211811 96 211827
rect 62 210819 96 210835
rect -50 210751 -34 210785
rect 34 210751 50 210785
rect -50 210643 -34 210677
rect 34 210643 50 210677
rect -96 210593 -62 210609
rect -96 209601 -62 209617
rect 62 210593 96 210609
rect 62 209601 96 209617
rect -50 209533 -34 209567
rect 34 209533 50 209567
rect -50 209425 -34 209459
rect 34 209425 50 209459
rect -96 209375 -62 209391
rect -96 208383 -62 208399
rect 62 209375 96 209391
rect 62 208383 96 208399
rect -50 208315 -34 208349
rect 34 208315 50 208349
rect -50 208207 -34 208241
rect 34 208207 50 208241
rect -96 208157 -62 208173
rect -96 207165 -62 207181
rect 62 208157 96 208173
rect 62 207165 96 207181
rect -50 207097 -34 207131
rect 34 207097 50 207131
rect -50 206989 -34 207023
rect 34 206989 50 207023
rect -96 206939 -62 206955
rect -96 205947 -62 205963
rect 62 206939 96 206955
rect 62 205947 96 205963
rect -50 205879 -34 205913
rect 34 205879 50 205913
rect -50 205771 -34 205805
rect 34 205771 50 205805
rect -96 205721 -62 205737
rect -96 204729 -62 204745
rect 62 205721 96 205737
rect 62 204729 96 204745
rect -50 204661 -34 204695
rect 34 204661 50 204695
rect -50 204553 -34 204587
rect 34 204553 50 204587
rect -96 204503 -62 204519
rect -96 203511 -62 203527
rect 62 204503 96 204519
rect 62 203511 96 203527
rect -50 203443 -34 203477
rect 34 203443 50 203477
rect -50 203335 -34 203369
rect 34 203335 50 203369
rect -96 203285 -62 203301
rect -96 202293 -62 202309
rect 62 203285 96 203301
rect 62 202293 96 202309
rect -50 202225 -34 202259
rect 34 202225 50 202259
rect -50 202117 -34 202151
rect 34 202117 50 202151
rect -96 202067 -62 202083
rect -96 201075 -62 201091
rect 62 202067 96 202083
rect 62 201075 96 201091
rect -50 201007 -34 201041
rect 34 201007 50 201041
rect -50 200899 -34 200933
rect 34 200899 50 200933
rect -96 200849 -62 200865
rect -96 199857 -62 199873
rect 62 200849 96 200865
rect 62 199857 96 199873
rect -50 199789 -34 199823
rect 34 199789 50 199823
rect -50 199681 -34 199715
rect 34 199681 50 199715
rect -96 199631 -62 199647
rect -96 198639 -62 198655
rect 62 199631 96 199647
rect 62 198639 96 198655
rect -50 198571 -34 198605
rect 34 198571 50 198605
rect -50 198463 -34 198497
rect 34 198463 50 198497
rect -96 198413 -62 198429
rect -96 197421 -62 197437
rect 62 198413 96 198429
rect 62 197421 96 197437
rect -50 197353 -34 197387
rect 34 197353 50 197387
rect -50 197245 -34 197279
rect 34 197245 50 197279
rect -96 197195 -62 197211
rect -96 196203 -62 196219
rect 62 197195 96 197211
rect 62 196203 96 196219
rect -50 196135 -34 196169
rect 34 196135 50 196169
rect -50 196027 -34 196061
rect 34 196027 50 196061
rect -96 195977 -62 195993
rect -96 194985 -62 195001
rect 62 195977 96 195993
rect 62 194985 96 195001
rect -50 194917 -34 194951
rect 34 194917 50 194951
rect -50 194809 -34 194843
rect 34 194809 50 194843
rect -96 194759 -62 194775
rect -96 193767 -62 193783
rect 62 194759 96 194775
rect 62 193767 96 193783
rect -50 193699 -34 193733
rect 34 193699 50 193733
rect -50 193591 -34 193625
rect 34 193591 50 193625
rect -96 193541 -62 193557
rect -96 192549 -62 192565
rect 62 193541 96 193557
rect 62 192549 96 192565
rect -50 192481 -34 192515
rect 34 192481 50 192515
rect -50 192373 -34 192407
rect 34 192373 50 192407
rect -96 192323 -62 192339
rect -96 191331 -62 191347
rect 62 192323 96 192339
rect 62 191331 96 191347
rect -50 191263 -34 191297
rect 34 191263 50 191297
rect -50 191155 -34 191189
rect 34 191155 50 191189
rect -96 191105 -62 191121
rect -96 190113 -62 190129
rect 62 191105 96 191121
rect 62 190113 96 190129
rect -50 190045 -34 190079
rect 34 190045 50 190079
rect -50 189937 -34 189971
rect 34 189937 50 189971
rect -96 189887 -62 189903
rect -96 188895 -62 188911
rect 62 189887 96 189903
rect 62 188895 96 188911
rect -50 188827 -34 188861
rect 34 188827 50 188861
rect -50 188719 -34 188753
rect 34 188719 50 188753
rect -96 188669 -62 188685
rect -96 187677 -62 187693
rect 62 188669 96 188685
rect 62 187677 96 187693
rect -50 187609 -34 187643
rect 34 187609 50 187643
rect -50 187501 -34 187535
rect 34 187501 50 187535
rect -96 187451 -62 187467
rect -96 186459 -62 186475
rect 62 187451 96 187467
rect 62 186459 96 186475
rect -50 186391 -34 186425
rect 34 186391 50 186425
rect -50 186283 -34 186317
rect 34 186283 50 186317
rect -96 186233 -62 186249
rect -96 185241 -62 185257
rect 62 186233 96 186249
rect 62 185241 96 185257
rect -50 185173 -34 185207
rect 34 185173 50 185207
rect -50 185065 -34 185099
rect 34 185065 50 185099
rect -96 185015 -62 185031
rect -96 184023 -62 184039
rect 62 185015 96 185031
rect 62 184023 96 184039
rect -50 183955 -34 183989
rect 34 183955 50 183989
rect -50 183847 -34 183881
rect 34 183847 50 183881
rect -96 183797 -62 183813
rect -96 182805 -62 182821
rect 62 183797 96 183813
rect 62 182805 96 182821
rect -50 182737 -34 182771
rect 34 182737 50 182771
rect -50 182629 -34 182663
rect 34 182629 50 182663
rect -96 182579 -62 182595
rect -96 181587 -62 181603
rect 62 182579 96 182595
rect 62 181587 96 181603
rect -50 181519 -34 181553
rect 34 181519 50 181553
rect -50 181411 -34 181445
rect 34 181411 50 181445
rect -96 181361 -62 181377
rect -96 180369 -62 180385
rect 62 181361 96 181377
rect 62 180369 96 180385
rect -50 180301 -34 180335
rect 34 180301 50 180335
rect -50 180193 -34 180227
rect 34 180193 50 180227
rect -96 180143 -62 180159
rect -96 179151 -62 179167
rect 62 180143 96 180159
rect 62 179151 96 179167
rect -50 179083 -34 179117
rect 34 179083 50 179117
rect -50 178975 -34 179009
rect 34 178975 50 179009
rect -96 178925 -62 178941
rect -96 177933 -62 177949
rect 62 178925 96 178941
rect 62 177933 96 177949
rect -50 177865 -34 177899
rect 34 177865 50 177899
rect -50 177757 -34 177791
rect 34 177757 50 177791
rect -96 177707 -62 177723
rect -96 176715 -62 176731
rect 62 177707 96 177723
rect 62 176715 96 176731
rect -50 176647 -34 176681
rect 34 176647 50 176681
rect -50 176539 -34 176573
rect 34 176539 50 176573
rect -96 176489 -62 176505
rect -96 175497 -62 175513
rect 62 176489 96 176505
rect 62 175497 96 175513
rect -50 175429 -34 175463
rect 34 175429 50 175463
rect -50 175321 -34 175355
rect 34 175321 50 175355
rect -96 175271 -62 175287
rect -96 174279 -62 174295
rect 62 175271 96 175287
rect 62 174279 96 174295
rect -50 174211 -34 174245
rect 34 174211 50 174245
rect -50 174103 -34 174137
rect 34 174103 50 174137
rect -96 174053 -62 174069
rect -96 173061 -62 173077
rect 62 174053 96 174069
rect 62 173061 96 173077
rect -50 172993 -34 173027
rect 34 172993 50 173027
rect -50 172885 -34 172919
rect 34 172885 50 172919
rect -96 172835 -62 172851
rect -96 171843 -62 171859
rect 62 172835 96 172851
rect 62 171843 96 171859
rect -50 171775 -34 171809
rect 34 171775 50 171809
rect -50 171667 -34 171701
rect 34 171667 50 171701
rect -96 171617 -62 171633
rect -96 170625 -62 170641
rect 62 171617 96 171633
rect 62 170625 96 170641
rect -50 170557 -34 170591
rect 34 170557 50 170591
rect -50 170449 -34 170483
rect 34 170449 50 170483
rect -96 170399 -62 170415
rect -96 169407 -62 169423
rect 62 170399 96 170415
rect 62 169407 96 169423
rect -50 169339 -34 169373
rect 34 169339 50 169373
rect -50 169231 -34 169265
rect 34 169231 50 169265
rect -96 169181 -62 169197
rect -96 168189 -62 168205
rect 62 169181 96 169197
rect 62 168189 96 168205
rect -50 168121 -34 168155
rect 34 168121 50 168155
rect -50 168013 -34 168047
rect 34 168013 50 168047
rect -96 167963 -62 167979
rect -96 166971 -62 166987
rect 62 167963 96 167979
rect 62 166971 96 166987
rect -50 166903 -34 166937
rect 34 166903 50 166937
rect -50 166795 -34 166829
rect 34 166795 50 166829
rect -96 166745 -62 166761
rect -96 165753 -62 165769
rect 62 166745 96 166761
rect 62 165753 96 165769
rect -50 165685 -34 165719
rect 34 165685 50 165719
rect -50 165577 -34 165611
rect 34 165577 50 165611
rect -96 165527 -62 165543
rect -96 164535 -62 164551
rect 62 165527 96 165543
rect 62 164535 96 164551
rect -50 164467 -34 164501
rect 34 164467 50 164501
rect -50 164359 -34 164393
rect 34 164359 50 164393
rect -96 164309 -62 164325
rect -96 163317 -62 163333
rect 62 164309 96 164325
rect 62 163317 96 163333
rect -50 163249 -34 163283
rect 34 163249 50 163283
rect -50 163141 -34 163175
rect 34 163141 50 163175
rect -96 163091 -62 163107
rect -96 162099 -62 162115
rect 62 163091 96 163107
rect 62 162099 96 162115
rect -50 162031 -34 162065
rect 34 162031 50 162065
rect -50 161923 -34 161957
rect 34 161923 50 161957
rect -96 161873 -62 161889
rect -96 160881 -62 160897
rect 62 161873 96 161889
rect 62 160881 96 160897
rect -50 160813 -34 160847
rect 34 160813 50 160847
rect -50 160705 -34 160739
rect 34 160705 50 160739
rect -96 160655 -62 160671
rect -96 159663 -62 159679
rect 62 160655 96 160671
rect 62 159663 96 159679
rect -50 159595 -34 159629
rect 34 159595 50 159629
rect -50 159487 -34 159521
rect 34 159487 50 159521
rect -96 159437 -62 159453
rect -96 158445 -62 158461
rect 62 159437 96 159453
rect 62 158445 96 158461
rect -50 158377 -34 158411
rect 34 158377 50 158411
rect -50 158269 -34 158303
rect 34 158269 50 158303
rect -96 158219 -62 158235
rect -96 157227 -62 157243
rect 62 158219 96 158235
rect 62 157227 96 157243
rect -50 157159 -34 157193
rect 34 157159 50 157193
rect -50 157051 -34 157085
rect 34 157051 50 157085
rect -96 157001 -62 157017
rect -96 156009 -62 156025
rect 62 157001 96 157017
rect 62 156009 96 156025
rect -50 155941 -34 155975
rect 34 155941 50 155975
rect -50 155833 -34 155867
rect 34 155833 50 155867
rect -96 155783 -62 155799
rect -96 154791 -62 154807
rect 62 155783 96 155799
rect 62 154791 96 154807
rect -50 154723 -34 154757
rect 34 154723 50 154757
rect -50 154615 -34 154649
rect 34 154615 50 154649
rect -96 154565 -62 154581
rect -96 153573 -62 153589
rect 62 154565 96 154581
rect 62 153573 96 153589
rect -50 153505 -34 153539
rect 34 153505 50 153539
rect -50 153397 -34 153431
rect 34 153397 50 153431
rect -96 153347 -62 153363
rect -96 152355 -62 152371
rect 62 153347 96 153363
rect 62 152355 96 152371
rect -50 152287 -34 152321
rect 34 152287 50 152321
rect -50 152179 -34 152213
rect 34 152179 50 152213
rect -96 152129 -62 152145
rect -96 151137 -62 151153
rect 62 152129 96 152145
rect 62 151137 96 151153
rect -50 151069 -34 151103
rect 34 151069 50 151103
rect -50 150961 -34 150995
rect 34 150961 50 150995
rect -96 150911 -62 150927
rect -96 149919 -62 149935
rect 62 150911 96 150927
rect 62 149919 96 149935
rect -50 149851 -34 149885
rect 34 149851 50 149885
rect -50 149743 -34 149777
rect 34 149743 50 149777
rect -96 149693 -62 149709
rect -96 148701 -62 148717
rect 62 149693 96 149709
rect 62 148701 96 148717
rect -50 148633 -34 148667
rect 34 148633 50 148667
rect -50 148525 -34 148559
rect 34 148525 50 148559
rect -96 148475 -62 148491
rect -96 147483 -62 147499
rect 62 148475 96 148491
rect 62 147483 96 147499
rect -50 147415 -34 147449
rect 34 147415 50 147449
rect -50 147307 -34 147341
rect 34 147307 50 147341
rect -96 147257 -62 147273
rect -96 146265 -62 146281
rect 62 147257 96 147273
rect 62 146265 96 146281
rect -50 146197 -34 146231
rect 34 146197 50 146231
rect -50 146089 -34 146123
rect 34 146089 50 146123
rect -96 146039 -62 146055
rect -96 145047 -62 145063
rect 62 146039 96 146055
rect 62 145047 96 145063
rect -50 144979 -34 145013
rect 34 144979 50 145013
rect -50 144871 -34 144905
rect 34 144871 50 144905
rect -96 144821 -62 144837
rect -96 143829 -62 143845
rect 62 144821 96 144837
rect 62 143829 96 143845
rect -50 143761 -34 143795
rect 34 143761 50 143795
rect -50 143653 -34 143687
rect 34 143653 50 143687
rect -96 143603 -62 143619
rect -96 142611 -62 142627
rect 62 143603 96 143619
rect 62 142611 96 142627
rect -50 142543 -34 142577
rect 34 142543 50 142577
rect -50 142435 -34 142469
rect 34 142435 50 142469
rect -96 142385 -62 142401
rect -96 141393 -62 141409
rect 62 142385 96 142401
rect 62 141393 96 141409
rect -50 141325 -34 141359
rect 34 141325 50 141359
rect -50 141217 -34 141251
rect 34 141217 50 141251
rect -96 141167 -62 141183
rect -96 140175 -62 140191
rect 62 141167 96 141183
rect 62 140175 96 140191
rect -50 140107 -34 140141
rect 34 140107 50 140141
rect -50 139999 -34 140033
rect 34 139999 50 140033
rect -96 139949 -62 139965
rect -96 138957 -62 138973
rect 62 139949 96 139965
rect 62 138957 96 138973
rect -50 138889 -34 138923
rect 34 138889 50 138923
rect -50 138781 -34 138815
rect 34 138781 50 138815
rect -96 138731 -62 138747
rect -96 137739 -62 137755
rect 62 138731 96 138747
rect 62 137739 96 137755
rect -50 137671 -34 137705
rect 34 137671 50 137705
rect -50 137563 -34 137597
rect 34 137563 50 137597
rect -96 137513 -62 137529
rect -96 136521 -62 136537
rect 62 137513 96 137529
rect 62 136521 96 136537
rect -50 136453 -34 136487
rect 34 136453 50 136487
rect -50 136345 -34 136379
rect 34 136345 50 136379
rect -96 136295 -62 136311
rect -96 135303 -62 135319
rect 62 136295 96 136311
rect 62 135303 96 135319
rect -50 135235 -34 135269
rect 34 135235 50 135269
rect -50 135127 -34 135161
rect 34 135127 50 135161
rect -96 135077 -62 135093
rect -96 134085 -62 134101
rect 62 135077 96 135093
rect 62 134085 96 134101
rect -50 134017 -34 134051
rect 34 134017 50 134051
rect -50 133909 -34 133943
rect 34 133909 50 133943
rect -96 133859 -62 133875
rect -96 132867 -62 132883
rect 62 133859 96 133875
rect 62 132867 96 132883
rect -50 132799 -34 132833
rect 34 132799 50 132833
rect -50 132691 -34 132725
rect 34 132691 50 132725
rect -96 132641 -62 132657
rect -96 131649 -62 131665
rect 62 132641 96 132657
rect 62 131649 96 131665
rect -50 131581 -34 131615
rect 34 131581 50 131615
rect -50 131473 -34 131507
rect 34 131473 50 131507
rect -96 131423 -62 131439
rect -96 130431 -62 130447
rect 62 131423 96 131439
rect 62 130431 96 130447
rect -50 130363 -34 130397
rect 34 130363 50 130397
rect -50 130255 -34 130289
rect 34 130255 50 130289
rect -96 130205 -62 130221
rect -96 129213 -62 129229
rect 62 130205 96 130221
rect 62 129213 96 129229
rect -50 129145 -34 129179
rect 34 129145 50 129179
rect -50 129037 -34 129071
rect 34 129037 50 129071
rect -96 128987 -62 129003
rect -96 127995 -62 128011
rect 62 128987 96 129003
rect 62 127995 96 128011
rect -50 127927 -34 127961
rect 34 127927 50 127961
rect -50 127819 -34 127853
rect 34 127819 50 127853
rect -96 127769 -62 127785
rect -96 126777 -62 126793
rect 62 127769 96 127785
rect 62 126777 96 126793
rect -50 126709 -34 126743
rect 34 126709 50 126743
rect -50 126601 -34 126635
rect 34 126601 50 126635
rect -96 126551 -62 126567
rect -96 125559 -62 125575
rect 62 126551 96 126567
rect 62 125559 96 125575
rect -50 125491 -34 125525
rect 34 125491 50 125525
rect -50 125383 -34 125417
rect 34 125383 50 125417
rect -96 125333 -62 125349
rect -96 124341 -62 124357
rect 62 125333 96 125349
rect 62 124341 96 124357
rect -50 124273 -34 124307
rect 34 124273 50 124307
rect -50 124165 -34 124199
rect 34 124165 50 124199
rect -96 124115 -62 124131
rect -96 123123 -62 123139
rect 62 124115 96 124131
rect 62 123123 96 123139
rect -50 123055 -34 123089
rect 34 123055 50 123089
rect -50 122947 -34 122981
rect 34 122947 50 122981
rect -96 122897 -62 122913
rect -96 121905 -62 121921
rect 62 122897 96 122913
rect 62 121905 96 121921
rect -50 121837 -34 121871
rect 34 121837 50 121871
rect -50 121729 -34 121763
rect 34 121729 50 121763
rect -96 121679 -62 121695
rect -96 120687 -62 120703
rect 62 121679 96 121695
rect 62 120687 96 120703
rect -50 120619 -34 120653
rect 34 120619 50 120653
rect -50 120511 -34 120545
rect 34 120511 50 120545
rect -96 120461 -62 120477
rect -96 119469 -62 119485
rect 62 120461 96 120477
rect 62 119469 96 119485
rect -50 119401 -34 119435
rect 34 119401 50 119435
rect -50 119293 -34 119327
rect 34 119293 50 119327
rect -96 119243 -62 119259
rect -96 118251 -62 118267
rect 62 119243 96 119259
rect 62 118251 96 118267
rect -50 118183 -34 118217
rect 34 118183 50 118217
rect -50 118075 -34 118109
rect 34 118075 50 118109
rect -96 118025 -62 118041
rect -96 117033 -62 117049
rect 62 118025 96 118041
rect 62 117033 96 117049
rect -50 116965 -34 116999
rect 34 116965 50 116999
rect -50 116857 -34 116891
rect 34 116857 50 116891
rect -96 116807 -62 116823
rect -96 115815 -62 115831
rect 62 116807 96 116823
rect 62 115815 96 115831
rect -50 115747 -34 115781
rect 34 115747 50 115781
rect -50 115639 -34 115673
rect 34 115639 50 115673
rect -96 115589 -62 115605
rect -96 114597 -62 114613
rect 62 115589 96 115605
rect 62 114597 96 114613
rect -50 114529 -34 114563
rect 34 114529 50 114563
rect -50 114421 -34 114455
rect 34 114421 50 114455
rect -96 114371 -62 114387
rect -96 113379 -62 113395
rect 62 114371 96 114387
rect 62 113379 96 113395
rect -50 113311 -34 113345
rect 34 113311 50 113345
rect -50 113203 -34 113237
rect 34 113203 50 113237
rect -96 113153 -62 113169
rect -96 112161 -62 112177
rect 62 113153 96 113169
rect 62 112161 96 112177
rect -50 112093 -34 112127
rect 34 112093 50 112127
rect -50 111985 -34 112019
rect 34 111985 50 112019
rect -96 111935 -62 111951
rect -96 110943 -62 110959
rect 62 111935 96 111951
rect 62 110943 96 110959
rect -50 110875 -34 110909
rect 34 110875 50 110909
rect -50 110767 -34 110801
rect 34 110767 50 110801
rect -96 110717 -62 110733
rect -96 109725 -62 109741
rect 62 110717 96 110733
rect 62 109725 96 109741
rect -50 109657 -34 109691
rect 34 109657 50 109691
rect -50 109549 -34 109583
rect 34 109549 50 109583
rect -96 109499 -62 109515
rect -96 108507 -62 108523
rect 62 109499 96 109515
rect 62 108507 96 108523
rect -50 108439 -34 108473
rect 34 108439 50 108473
rect -50 108331 -34 108365
rect 34 108331 50 108365
rect -96 108281 -62 108297
rect -96 107289 -62 107305
rect 62 108281 96 108297
rect 62 107289 96 107305
rect -50 107221 -34 107255
rect 34 107221 50 107255
rect -50 107113 -34 107147
rect 34 107113 50 107147
rect -96 107063 -62 107079
rect -96 106071 -62 106087
rect 62 107063 96 107079
rect 62 106071 96 106087
rect -50 106003 -34 106037
rect 34 106003 50 106037
rect -50 105895 -34 105929
rect 34 105895 50 105929
rect -96 105845 -62 105861
rect -96 104853 -62 104869
rect 62 105845 96 105861
rect 62 104853 96 104869
rect -50 104785 -34 104819
rect 34 104785 50 104819
rect -50 104677 -34 104711
rect 34 104677 50 104711
rect -96 104627 -62 104643
rect -96 103635 -62 103651
rect 62 104627 96 104643
rect 62 103635 96 103651
rect -50 103567 -34 103601
rect 34 103567 50 103601
rect -50 103459 -34 103493
rect 34 103459 50 103493
rect -96 103409 -62 103425
rect -96 102417 -62 102433
rect 62 103409 96 103425
rect 62 102417 96 102433
rect -50 102349 -34 102383
rect 34 102349 50 102383
rect -50 102241 -34 102275
rect 34 102241 50 102275
rect -96 102191 -62 102207
rect -96 101199 -62 101215
rect 62 102191 96 102207
rect 62 101199 96 101215
rect -50 101131 -34 101165
rect 34 101131 50 101165
rect -50 101023 -34 101057
rect 34 101023 50 101057
rect -96 100973 -62 100989
rect -96 99981 -62 99997
rect 62 100973 96 100989
rect 62 99981 96 99997
rect -50 99913 -34 99947
rect 34 99913 50 99947
rect -50 99805 -34 99839
rect 34 99805 50 99839
rect -96 99755 -62 99771
rect -96 98763 -62 98779
rect 62 99755 96 99771
rect 62 98763 96 98779
rect -50 98695 -34 98729
rect 34 98695 50 98729
rect -50 98587 -34 98621
rect 34 98587 50 98621
rect -96 98537 -62 98553
rect -96 97545 -62 97561
rect 62 98537 96 98553
rect 62 97545 96 97561
rect -50 97477 -34 97511
rect 34 97477 50 97511
rect -50 97369 -34 97403
rect 34 97369 50 97403
rect -96 97319 -62 97335
rect -96 96327 -62 96343
rect 62 97319 96 97335
rect 62 96327 96 96343
rect -50 96259 -34 96293
rect 34 96259 50 96293
rect -50 96151 -34 96185
rect 34 96151 50 96185
rect -96 96101 -62 96117
rect -96 95109 -62 95125
rect 62 96101 96 96117
rect 62 95109 96 95125
rect -50 95041 -34 95075
rect 34 95041 50 95075
rect -50 94933 -34 94967
rect 34 94933 50 94967
rect -96 94883 -62 94899
rect -96 93891 -62 93907
rect 62 94883 96 94899
rect 62 93891 96 93907
rect -50 93823 -34 93857
rect 34 93823 50 93857
rect -50 93715 -34 93749
rect 34 93715 50 93749
rect -96 93665 -62 93681
rect -96 92673 -62 92689
rect 62 93665 96 93681
rect 62 92673 96 92689
rect -50 92605 -34 92639
rect 34 92605 50 92639
rect -50 92497 -34 92531
rect 34 92497 50 92531
rect -96 92447 -62 92463
rect -96 91455 -62 91471
rect 62 92447 96 92463
rect 62 91455 96 91471
rect -50 91387 -34 91421
rect 34 91387 50 91421
rect -50 91279 -34 91313
rect 34 91279 50 91313
rect -96 91229 -62 91245
rect -96 90237 -62 90253
rect 62 91229 96 91245
rect 62 90237 96 90253
rect -50 90169 -34 90203
rect 34 90169 50 90203
rect -50 90061 -34 90095
rect 34 90061 50 90095
rect -96 90011 -62 90027
rect -96 89019 -62 89035
rect 62 90011 96 90027
rect 62 89019 96 89035
rect -50 88951 -34 88985
rect 34 88951 50 88985
rect -50 88843 -34 88877
rect 34 88843 50 88877
rect -96 88793 -62 88809
rect -96 87801 -62 87817
rect 62 88793 96 88809
rect 62 87801 96 87817
rect -50 87733 -34 87767
rect 34 87733 50 87767
rect -50 87625 -34 87659
rect 34 87625 50 87659
rect -96 87575 -62 87591
rect -96 86583 -62 86599
rect 62 87575 96 87591
rect 62 86583 96 86599
rect -50 86515 -34 86549
rect 34 86515 50 86549
rect -50 86407 -34 86441
rect 34 86407 50 86441
rect -96 86357 -62 86373
rect -96 85365 -62 85381
rect 62 86357 96 86373
rect 62 85365 96 85381
rect -50 85297 -34 85331
rect 34 85297 50 85331
rect -50 85189 -34 85223
rect 34 85189 50 85223
rect -96 85139 -62 85155
rect -96 84147 -62 84163
rect 62 85139 96 85155
rect 62 84147 96 84163
rect -50 84079 -34 84113
rect 34 84079 50 84113
rect -50 83971 -34 84005
rect 34 83971 50 84005
rect -96 83921 -62 83937
rect -96 82929 -62 82945
rect 62 83921 96 83937
rect 62 82929 96 82945
rect -50 82861 -34 82895
rect 34 82861 50 82895
rect -50 82753 -34 82787
rect 34 82753 50 82787
rect -96 82703 -62 82719
rect -96 81711 -62 81727
rect 62 82703 96 82719
rect 62 81711 96 81727
rect -50 81643 -34 81677
rect 34 81643 50 81677
rect -50 81535 -34 81569
rect 34 81535 50 81569
rect -96 81485 -62 81501
rect -96 80493 -62 80509
rect 62 81485 96 81501
rect 62 80493 96 80509
rect -50 80425 -34 80459
rect 34 80425 50 80459
rect -50 80317 -34 80351
rect 34 80317 50 80351
rect -96 80267 -62 80283
rect -96 79275 -62 79291
rect 62 80267 96 80283
rect 62 79275 96 79291
rect -50 79207 -34 79241
rect 34 79207 50 79241
rect -50 79099 -34 79133
rect 34 79099 50 79133
rect -96 79049 -62 79065
rect -96 78057 -62 78073
rect 62 79049 96 79065
rect 62 78057 96 78073
rect -50 77989 -34 78023
rect 34 77989 50 78023
rect -50 77881 -34 77915
rect 34 77881 50 77915
rect -96 77831 -62 77847
rect -96 76839 -62 76855
rect 62 77831 96 77847
rect 62 76839 96 76855
rect -50 76771 -34 76805
rect 34 76771 50 76805
rect -50 76663 -34 76697
rect 34 76663 50 76697
rect -96 76613 -62 76629
rect -96 75621 -62 75637
rect 62 76613 96 76629
rect 62 75621 96 75637
rect -50 75553 -34 75587
rect 34 75553 50 75587
rect -50 75445 -34 75479
rect 34 75445 50 75479
rect -96 75395 -62 75411
rect -96 74403 -62 74419
rect 62 75395 96 75411
rect 62 74403 96 74419
rect -50 74335 -34 74369
rect 34 74335 50 74369
rect -50 74227 -34 74261
rect 34 74227 50 74261
rect -96 74177 -62 74193
rect -96 73185 -62 73201
rect 62 74177 96 74193
rect 62 73185 96 73201
rect -50 73117 -34 73151
rect 34 73117 50 73151
rect -50 73009 -34 73043
rect 34 73009 50 73043
rect -96 72959 -62 72975
rect -96 71967 -62 71983
rect 62 72959 96 72975
rect 62 71967 96 71983
rect -50 71899 -34 71933
rect 34 71899 50 71933
rect -50 71791 -34 71825
rect 34 71791 50 71825
rect -96 71741 -62 71757
rect -96 70749 -62 70765
rect 62 71741 96 71757
rect 62 70749 96 70765
rect -50 70681 -34 70715
rect 34 70681 50 70715
rect -50 70573 -34 70607
rect 34 70573 50 70607
rect -96 70523 -62 70539
rect -96 69531 -62 69547
rect 62 70523 96 70539
rect 62 69531 96 69547
rect -50 69463 -34 69497
rect 34 69463 50 69497
rect -50 69355 -34 69389
rect 34 69355 50 69389
rect -96 69305 -62 69321
rect -96 68313 -62 68329
rect 62 69305 96 69321
rect 62 68313 96 68329
rect -50 68245 -34 68279
rect 34 68245 50 68279
rect -50 68137 -34 68171
rect 34 68137 50 68171
rect -96 68087 -62 68103
rect -96 67095 -62 67111
rect 62 68087 96 68103
rect 62 67095 96 67111
rect -50 67027 -34 67061
rect 34 67027 50 67061
rect -50 66919 -34 66953
rect 34 66919 50 66953
rect -96 66869 -62 66885
rect -96 65877 -62 65893
rect 62 66869 96 66885
rect 62 65877 96 65893
rect -50 65809 -34 65843
rect 34 65809 50 65843
rect -50 65701 -34 65735
rect 34 65701 50 65735
rect -96 65651 -62 65667
rect -96 64659 -62 64675
rect 62 65651 96 65667
rect 62 64659 96 64675
rect -50 64591 -34 64625
rect 34 64591 50 64625
rect -50 64483 -34 64517
rect 34 64483 50 64517
rect -96 64433 -62 64449
rect -96 63441 -62 63457
rect 62 64433 96 64449
rect 62 63441 96 63457
rect -50 63373 -34 63407
rect 34 63373 50 63407
rect -50 63265 -34 63299
rect 34 63265 50 63299
rect -96 63215 -62 63231
rect -96 62223 -62 62239
rect 62 63215 96 63231
rect 62 62223 96 62239
rect -50 62155 -34 62189
rect 34 62155 50 62189
rect -50 62047 -34 62081
rect 34 62047 50 62081
rect -96 61997 -62 62013
rect -96 61005 -62 61021
rect 62 61997 96 62013
rect 62 61005 96 61021
rect -50 60937 -34 60971
rect 34 60937 50 60971
rect -50 60829 -34 60863
rect 34 60829 50 60863
rect -96 60779 -62 60795
rect -96 59787 -62 59803
rect 62 60779 96 60795
rect 62 59787 96 59803
rect -50 59719 -34 59753
rect 34 59719 50 59753
rect -50 59611 -34 59645
rect 34 59611 50 59645
rect -96 59561 -62 59577
rect -96 58569 -62 58585
rect 62 59561 96 59577
rect 62 58569 96 58585
rect -50 58501 -34 58535
rect 34 58501 50 58535
rect -50 58393 -34 58427
rect 34 58393 50 58427
rect -96 58343 -62 58359
rect -96 57351 -62 57367
rect 62 58343 96 58359
rect 62 57351 96 57367
rect -50 57283 -34 57317
rect 34 57283 50 57317
rect -50 57175 -34 57209
rect 34 57175 50 57209
rect -96 57125 -62 57141
rect -96 56133 -62 56149
rect 62 57125 96 57141
rect 62 56133 96 56149
rect -50 56065 -34 56099
rect 34 56065 50 56099
rect -50 55957 -34 55991
rect 34 55957 50 55991
rect -96 55907 -62 55923
rect -96 54915 -62 54931
rect 62 55907 96 55923
rect 62 54915 96 54931
rect -50 54847 -34 54881
rect 34 54847 50 54881
rect -50 54739 -34 54773
rect 34 54739 50 54773
rect -96 54689 -62 54705
rect -96 53697 -62 53713
rect 62 54689 96 54705
rect 62 53697 96 53713
rect -50 53629 -34 53663
rect 34 53629 50 53663
rect -50 53521 -34 53555
rect 34 53521 50 53555
rect -96 53471 -62 53487
rect -96 52479 -62 52495
rect 62 53471 96 53487
rect 62 52479 96 52495
rect -50 52411 -34 52445
rect 34 52411 50 52445
rect -50 52303 -34 52337
rect 34 52303 50 52337
rect -96 52253 -62 52269
rect -96 51261 -62 51277
rect 62 52253 96 52269
rect 62 51261 96 51277
rect -50 51193 -34 51227
rect 34 51193 50 51227
rect -50 51085 -34 51119
rect 34 51085 50 51119
rect -96 51035 -62 51051
rect -96 50043 -62 50059
rect 62 51035 96 51051
rect 62 50043 96 50059
rect -50 49975 -34 50009
rect 34 49975 50 50009
rect -50 49867 -34 49901
rect 34 49867 50 49901
rect -96 49817 -62 49833
rect -96 48825 -62 48841
rect 62 49817 96 49833
rect 62 48825 96 48841
rect -50 48757 -34 48791
rect 34 48757 50 48791
rect -50 48649 -34 48683
rect 34 48649 50 48683
rect -96 48599 -62 48615
rect -96 47607 -62 47623
rect 62 48599 96 48615
rect 62 47607 96 47623
rect -50 47539 -34 47573
rect 34 47539 50 47573
rect -50 47431 -34 47465
rect 34 47431 50 47465
rect -96 47381 -62 47397
rect -96 46389 -62 46405
rect 62 47381 96 47397
rect 62 46389 96 46405
rect -50 46321 -34 46355
rect 34 46321 50 46355
rect -50 46213 -34 46247
rect 34 46213 50 46247
rect -96 46163 -62 46179
rect -96 45171 -62 45187
rect 62 46163 96 46179
rect 62 45171 96 45187
rect -50 45103 -34 45137
rect 34 45103 50 45137
rect -50 44995 -34 45029
rect 34 44995 50 45029
rect -96 44945 -62 44961
rect -96 43953 -62 43969
rect 62 44945 96 44961
rect 62 43953 96 43969
rect -50 43885 -34 43919
rect 34 43885 50 43919
rect -50 43777 -34 43811
rect 34 43777 50 43811
rect -96 43727 -62 43743
rect -96 42735 -62 42751
rect 62 43727 96 43743
rect 62 42735 96 42751
rect -50 42667 -34 42701
rect 34 42667 50 42701
rect -50 42559 -34 42593
rect 34 42559 50 42593
rect -96 42509 -62 42525
rect -96 41517 -62 41533
rect 62 42509 96 42525
rect 62 41517 96 41533
rect -50 41449 -34 41483
rect 34 41449 50 41483
rect -50 41341 -34 41375
rect 34 41341 50 41375
rect -96 41291 -62 41307
rect -96 40299 -62 40315
rect 62 41291 96 41307
rect 62 40299 96 40315
rect -50 40231 -34 40265
rect 34 40231 50 40265
rect -50 40123 -34 40157
rect 34 40123 50 40157
rect -96 40073 -62 40089
rect -96 39081 -62 39097
rect 62 40073 96 40089
rect 62 39081 96 39097
rect -50 39013 -34 39047
rect 34 39013 50 39047
rect -50 38905 -34 38939
rect 34 38905 50 38939
rect -96 38855 -62 38871
rect -96 37863 -62 37879
rect 62 38855 96 38871
rect 62 37863 96 37879
rect -50 37795 -34 37829
rect 34 37795 50 37829
rect -50 37687 -34 37721
rect 34 37687 50 37721
rect -96 37637 -62 37653
rect -96 36645 -62 36661
rect 62 37637 96 37653
rect 62 36645 96 36661
rect -50 36577 -34 36611
rect 34 36577 50 36611
rect -50 36469 -34 36503
rect 34 36469 50 36503
rect -96 36419 -62 36435
rect -96 35427 -62 35443
rect 62 36419 96 36435
rect 62 35427 96 35443
rect -50 35359 -34 35393
rect 34 35359 50 35393
rect -50 35251 -34 35285
rect 34 35251 50 35285
rect -96 35201 -62 35217
rect -96 34209 -62 34225
rect 62 35201 96 35217
rect 62 34209 96 34225
rect -50 34141 -34 34175
rect 34 34141 50 34175
rect -50 34033 -34 34067
rect 34 34033 50 34067
rect -96 33983 -62 33999
rect -96 32991 -62 33007
rect 62 33983 96 33999
rect 62 32991 96 33007
rect -50 32923 -34 32957
rect 34 32923 50 32957
rect -50 32815 -34 32849
rect 34 32815 50 32849
rect -96 32765 -62 32781
rect -96 31773 -62 31789
rect 62 32765 96 32781
rect 62 31773 96 31789
rect -50 31705 -34 31739
rect 34 31705 50 31739
rect -50 31597 -34 31631
rect 34 31597 50 31631
rect -96 31547 -62 31563
rect -96 30555 -62 30571
rect 62 31547 96 31563
rect 62 30555 96 30571
rect -50 30487 -34 30521
rect 34 30487 50 30521
rect -50 30379 -34 30413
rect 34 30379 50 30413
rect -96 30329 -62 30345
rect -96 29337 -62 29353
rect 62 30329 96 30345
rect 62 29337 96 29353
rect -50 29269 -34 29303
rect 34 29269 50 29303
rect -50 29161 -34 29195
rect 34 29161 50 29195
rect -96 29111 -62 29127
rect -96 28119 -62 28135
rect 62 29111 96 29127
rect 62 28119 96 28135
rect -50 28051 -34 28085
rect 34 28051 50 28085
rect -50 27943 -34 27977
rect 34 27943 50 27977
rect -96 27893 -62 27909
rect -96 26901 -62 26917
rect 62 27893 96 27909
rect 62 26901 96 26917
rect -50 26833 -34 26867
rect 34 26833 50 26867
rect -50 26725 -34 26759
rect 34 26725 50 26759
rect -96 26675 -62 26691
rect -96 25683 -62 25699
rect 62 26675 96 26691
rect 62 25683 96 25699
rect -50 25615 -34 25649
rect 34 25615 50 25649
rect -50 25507 -34 25541
rect 34 25507 50 25541
rect -96 25457 -62 25473
rect -96 24465 -62 24481
rect 62 25457 96 25473
rect 62 24465 96 24481
rect -50 24397 -34 24431
rect 34 24397 50 24431
rect -50 24289 -34 24323
rect 34 24289 50 24323
rect -96 24239 -62 24255
rect -96 23247 -62 23263
rect 62 24239 96 24255
rect 62 23247 96 23263
rect -50 23179 -34 23213
rect 34 23179 50 23213
rect -50 23071 -34 23105
rect 34 23071 50 23105
rect -96 23021 -62 23037
rect -96 22029 -62 22045
rect 62 23021 96 23037
rect 62 22029 96 22045
rect -50 21961 -34 21995
rect 34 21961 50 21995
rect -50 21853 -34 21887
rect 34 21853 50 21887
rect -96 21803 -62 21819
rect -96 20811 -62 20827
rect 62 21803 96 21819
rect 62 20811 96 20827
rect -50 20743 -34 20777
rect 34 20743 50 20777
rect -50 20635 -34 20669
rect 34 20635 50 20669
rect -96 20585 -62 20601
rect -96 19593 -62 19609
rect 62 20585 96 20601
rect 62 19593 96 19609
rect -50 19525 -34 19559
rect 34 19525 50 19559
rect -50 19417 -34 19451
rect 34 19417 50 19451
rect -96 19367 -62 19383
rect -96 18375 -62 18391
rect 62 19367 96 19383
rect 62 18375 96 18391
rect -50 18307 -34 18341
rect 34 18307 50 18341
rect -50 18199 -34 18233
rect 34 18199 50 18233
rect -96 18149 -62 18165
rect -96 17157 -62 17173
rect 62 18149 96 18165
rect 62 17157 96 17173
rect -50 17089 -34 17123
rect 34 17089 50 17123
rect -50 16981 -34 17015
rect 34 16981 50 17015
rect -96 16931 -62 16947
rect -96 15939 -62 15955
rect 62 16931 96 16947
rect 62 15939 96 15955
rect -50 15871 -34 15905
rect 34 15871 50 15905
rect -50 15763 -34 15797
rect 34 15763 50 15797
rect -96 15713 -62 15729
rect -96 14721 -62 14737
rect 62 15713 96 15729
rect 62 14721 96 14737
rect -50 14653 -34 14687
rect 34 14653 50 14687
rect -50 14545 -34 14579
rect 34 14545 50 14579
rect -96 14495 -62 14511
rect -96 13503 -62 13519
rect 62 14495 96 14511
rect 62 13503 96 13519
rect -50 13435 -34 13469
rect 34 13435 50 13469
rect -50 13327 -34 13361
rect 34 13327 50 13361
rect -96 13277 -62 13293
rect -96 12285 -62 12301
rect 62 13277 96 13293
rect 62 12285 96 12301
rect -50 12217 -34 12251
rect 34 12217 50 12251
rect -50 12109 -34 12143
rect 34 12109 50 12143
rect -96 12059 -62 12075
rect -96 11067 -62 11083
rect 62 12059 96 12075
rect 62 11067 96 11083
rect -50 10999 -34 11033
rect 34 10999 50 11033
rect -50 10891 -34 10925
rect 34 10891 50 10925
rect -96 10841 -62 10857
rect -96 9849 -62 9865
rect 62 10841 96 10857
rect 62 9849 96 9865
rect -50 9781 -34 9815
rect 34 9781 50 9815
rect -50 9673 -34 9707
rect 34 9673 50 9707
rect -96 9623 -62 9639
rect -96 8631 -62 8647
rect 62 9623 96 9639
rect 62 8631 96 8647
rect -50 8563 -34 8597
rect 34 8563 50 8597
rect -50 8455 -34 8489
rect 34 8455 50 8489
rect -96 8405 -62 8421
rect -96 7413 -62 7429
rect 62 8405 96 8421
rect 62 7413 96 7429
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -50 7237 -34 7271
rect 34 7237 50 7271
rect -96 7187 -62 7203
rect -96 6195 -62 6211
rect 62 7187 96 7203
rect 62 6195 96 6211
rect -50 6127 -34 6161
rect 34 6127 50 6161
rect -50 6019 -34 6053
rect 34 6019 50 6053
rect -96 5969 -62 5985
rect -96 4977 -62 4993
rect 62 5969 96 5985
rect 62 4977 96 4993
rect -50 4909 -34 4943
rect 34 4909 50 4943
rect -50 4801 -34 4835
rect 34 4801 50 4835
rect -96 4751 -62 4767
rect -96 3759 -62 3775
rect 62 4751 96 4767
rect 62 3759 96 3775
rect -50 3691 -34 3725
rect 34 3691 50 3725
rect -50 3583 -34 3617
rect 34 3583 50 3617
rect -96 3533 -62 3549
rect -96 2541 -62 2557
rect 62 3533 96 3549
rect 62 2541 96 2557
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -96 2315 -62 2331
rect -96 1323 -62 1339
rect 62 2315 96 2331
rect 62 1323 96 1339
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -96 1097 -62 1113
rect -96 105 -62 121
rect 62 1097 96 1113
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -1113 -62 -1097
rect 62 -121 96 -105
rect 62 -1113 96 -1097
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -96 -1339 -62 -1323
rect -96 -2331 -62 -2315
rect 62 -1339 96 -1323
rect 62 -2331 96 -2315
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -96 -2557 -62 -2541
rect -96 -3549 -62 -3533
rect 62 -2557 96 -2541
rect 62 -3549 96 -3533
rect -50 -3617 -34 -3583
rect 34 -3617 50 -3583
rect -50 -3725 -34 -3691
rect 34 -3725 50 -3691
rect -96 -3775 -62 -3759
rect -96 -4767 -62 -4751
rect 62 -3775 96 -3759
rect 62 -4767 96 -4751
rect -50 -4835 -34 -4801
rect 34 -4835 50 -4801
rect -50 -4943 -34 -4909
rect 34 -4943 50 -4909
rect -96 -4993 -62 -4977
rect -96 -5985 -62 -5969
rect 62 -4993 96 -4977
rect 62 -5985 96 -5969
rect -50 -6053 -34 -6019
rect 34 -6053 50 -6019
rect -50 -6161 -34 -6127
rect 34 -6161 50 -6127
rect -96 -6211 -62 -6195
rect -96 -7203 -62 -7187
rect 62 -6211 96 -6195
rect 62 -7203 96 -7187
rect -50 -7271 -34 -7237
rect 34 -7271 50 -7237
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -96 -7429 -62 -7413
rect -96 -8421 -62 -8405
rect 62 -7429 96 -7413
rect 62 -8421 96 -8405
rect -50 -8489 -34 -8455
rect 34 -8489 50 -8455
rect -50 -8597 -34 -8563
rect 34 -8597 50 -8563
rect -96 -8647 -62 -8631
rect -96 -9639 -62 -9623
rect 62 -8647 96 -8631
rect 62 -9639 96 -9623
rect -50 -9707 -34 -9673
rect 34 -9707 50 -9673
rect -50 -9815 -34 -9781
rect 34 -9815 50 -9781
rect -96 -9865 -62 -9849
rect -96 -10857 -62 -10841
rect 62 -9865 96 -9849
rect 62 -10857 96 -10841
rect -50 -10925 -34 -10891
rect 34 -10925 50 -10891
rect -50 -11033 -34 -10999
rect 34 -11033 50 -10999
rect -96 -11083 -62 -11067
rect -96 -12075 -62 -12059
rect 62 -11083 96 -11067
rect 62 -12075 96 -12059
rect -50 -12143 -34 -12109
rect 34 -12143 50 -12109
rect -50 -12251 -34 -12217
rect 34 -12251 50 -12217
rect -96 -12301 -62 -12285
rect -96 -13293 -62 -13277
rect 62 -12301 96 -12285
rect 62 -13293 96 -13277
rect -50 -13361 -34 -13327
rect 34 -13361 50 -13327
rect -50 -13469 -34 -13435
rect 34 -13469 50 -13435
rect -96 -13519 -62 -13503
rect -96 -14511 -62 -14495
rect 62 -13519 96 -13503
rect 62 -14511 96 -14495
rect -50 -14579 -34 -14545
rect 34 -14579 50 -14545
rect -50 -14687 -34 -14653
rect 34 -14687 50 -14653
rect -96 -14737 -62 -14721
rect -96 -15729 -62 -15713
rect 62 -14737 96 -14721
rect 62 -15729 96 -15713
rect -50 -15797 -34 -15763
rect 34 -15797 50 -15763
rect -50 -15905 -34 -15871
rect 34 -15905 50 -15871
rect -96 -15955 -62 -15939
rect -96 -16947 -62 -16931
rect 62 -15955 96 -15939
rect 62 -16947 96 -16931
rect -50 -17015 -34 -16981
rect 34 -17015 50 -16981
rect -50 -17123 -34 -17089
rect 34 -17123 50 -17089
rect -96 -17173 -62 -17157
rect -96 -18165 -62 -18149
rect 62 -17173 96 -17157
rect 62 -18165 96 -18149
rect -50 -18233 -34 -18199
rect 34 -18233 50 -18199
rect -50 -18341 -34 -18307
rect 34 -18341 50 -18307
rect -96 -18391 -62 -18375
rect -96 -19383 -62 -19367
rect 62 -18391 96 -18375
rect 62 -19383 96 -19367
rect -50 -19451 -34 -19417
rect 34 -19451 50 -19417
rect -50 -19559 -34 -19525
rect 34 -19559 50 -19525
rect -96 -19609 -62 -19593
rect -96 -20601 -62 -20585
rect 62 -19609 96 -19593
rect 62 -20601 96 -20585
rect -50 -20669 -34 -20635
rect 34 -20669 50 -20635
rect -50 -20777 -34 -20743
rect 34 -20777 50 -20743
rect -96 -20827 -62 -20811
rect -96 -21819 -62 -21803
rect 62 -20827 96 -20811
rect 62 -21819 96 -21803
rect -50 -21887 -34 -21853
rect 34 -21887 50 -21853
rect -50 -21995 -34 -21961
rect 34 -21995 50 -21961
rect -96 -22045 -62 -22029
rect -96 -23037 -62 -23021
rect 62 -22045 96 -22029
rect 62 -23037 96 -23021
rect -50 -23105 -34 -23071
rect 34 -23105 50 -23071
rect -50 -23213 -34 -23179
rect 34 -23213 50 -23179
rect -96 -23263 -62 -23247
rect -96 -24255 -62 -24239
rect 62 -23263 96 -23247
rect 62 -24255 96 -24239
rect -50 -24323 -34 -24289
rect 34 -24323 50 -24289
rect -50 -24431 -34 -24397
rect 34 -24431 50 -24397
rect -96 -24481 -62 -24465
rect -96 -25473 -62 -25457
rect 62 -24481 96 -24465
rect 62 -25473 96 -25457
rect -50 -25541 -34 -25507
rect 34 -25541 50 -25507
rect -50 -25649 -34 -25615
rect 34 -25649 50 -25615
rect -96 -25699 -62 -25683
rect -96 -26691 -62 -26675
rect 62 -25699 96 -25683
rect 62 -26691 96 -26675
rect -50 -26759 -34 -26725
rect 34 -26759 50 -26725
rect -50 -26867 -34 -26833
rect 34 -26867 50 -26833
rect -96 -26917 -62 -26901
rect -96 -27909 -62 -27893
rect 62 -26917 96 -26901
rect 62 -27909 96 -27893
rect -50 -27977 -34 -27943
rect 34 -27977 50 -27943
rect -50 -28085 -34 -28051
rect 34 -28085 50 -28051
rect -96 -28135 -62 -28119
rect -96 -29127 -62 -29111
rect 62 -28135 96 -28119
rect 62 -29127 96 -29111
rect -50 -29195 -34 -29161
rect 34 -29195 50 -29161
rect -50 -29303 -34 -29269
rect 34 -29303 50 -29269
rect -96 -29353 -62 -29337
rect -96 -30345 -62 -30329
rect 62 -29353 96 -29337
rect 62 -30345 96 -30329
rect -50 -30413 -34 -30379
rect 34 -30413 50 -30379
rect -50 -30521 -34 -30487
rect 34 -30521 50 -30487
rect -96 -30571 -62 -30555
rect -96 -31563 -62 -31547
rect 62 -30571 96 -30555
rect 62 -31563 96 -31547
rect -50 -31631 -34 -31597
rect 34 -31631 50 -31597
rect -50 -31739 -34 -31705
rect 34 -31739 50 -31705
rect -96 -31789 -62 -31773
rect -96 -32781 -62 -32765
rect 62 -31789 96 -31773
rect 62 -32781 96 -32765
rect -50 -32849 -34 -32815
rect 34 -32849 50 -32815
rect -50 -32957 -34 -32923
rect 34 -32957 50 -32923
rect -96 -33007 -62 -32991
rect -96 -33999 -62 -33983
rect 62 -33007 96 -32991
rect 62 -33999 96 -33983
rect -50 -34067 -34 -34033
rect 34 -34067 50 -34033
rect -50 -34175 -34 -34141
rect 34 -34175 50 -34141
rect -96 -34225 -62 -34209
rect -96 -35217 -62 -35201
rect 62 -34225 96 -34209
rect 62 -35217 96 -35201
rect -50 -35285 -34 -35251
rect 34 -35285 50 -35251
rect -50 -35393 -34 -35359
rect 34 -35393 50 -35359
rect -96 -35443 -62 -35427
rect -96 -36435 -62 -36419
rect 62 -35443 96 -35427
rect 62 -36435 96 -36419
rect -50 -36503 -34 -36469
rect 34 -36503 50 -36469
rect -50 -36611 -34 -36577
rect 34 -36611 50 -36577
rect -96 -36661 -62 -36645
rect -96 -37653 -62 -37637
rect 62 -36661 96 -36645
rect 62 -37653 96 -37637
rect -50 -37721 -34 -37687
rect 34 -37721 50 -37687
rect -50 -37829 -34 -37795
rect 34 -37829 50 -37795
rect -96 -37879 -62 -37863
rect -96 -38871 -62 -38855
rect 62 -37879 96 -37863
rect 62 -38871 96 -38855
rect -50 -38939 -34 -38905
rect 34 -38939 50 -38905
rect -50 -39047 -34 -39013
rect 34 -39047 50 -39013
rect -96 -39097 -62 -39081
rect -96 -40089 -62 -40073
rect 62 -39097 96 -39081
rect 62 -40089 96 -40073
rect -50 -40157 -34 -40123
rect 34 -40157 50 -40123
rect -50 -40265 -34 -40231
rect 34 -40265 50 -40231
rect -96 -40315 -62 -40299
rect -96 -41307 -62 -41291
rect 62 -40315 96 -40299
rect 62 -41307 96 -41291
rect -50 -41375 -34 -41341
rect 34 -41375 50 -41341
rect -50 -41483 -34 -41449
rect 34 -41483 50 -41449
rect -96 -41533 -62 -41517
rect -96 -42525 -62 -42509
rect 62 -41533 96 -41517
rect 62 -42525 96 -42509
rect -50 -42593 -34 -42559
rect 34 -42593 50 -42559
rect -50 -42701 -34 -42667
rect 34 -42701 50 -42667
rect -96 -42751 -62 -42735
rect -96 -43743 -62 -43727
rect 62 -42751 96 -42735
rect 62 -43743 96 -43727
rect -50 -43811 -34 -43777
rect 34 -43811 50 -43777
rect -50 -43919 -34 -43885
rect 34 -43919 50 -43885
rect -96 -43969 -62 -43953
rect -96 -44961 -62 -44945
rect 62 -43969 96 -43953
rect 62 -44961 96 -44945
rect -50 -45029 -34 -44995
rect 34 -45029 50 -44995
rect -50 -45137 -34 -45103
rect 34 -45137 50 -45103
rect -96 -45187 -62 -45171
rect -96 -46179 -62 -46163
rect 62 -45187 96 -45171
rect 62 -46179 96 -46163
rect -50 -46247 -34 -46213
rect 34 -46247 50 -46213
rect -50 -46355 -34 -46321
rect 34 -46355 50 -46321
rect -96 -46405 -62 -46389
rect -96 -47397 -62 -47381
rect 62 -46405 96 -46389
rect 62 -47397 96 -47381
rect -50 -47465 -34 -47431
rect 34 -47465 50 -47431
rect -50 -47573 -34 -47539
rect 34 -47573 50 -47539
rect -96 -47623 -62 -47607
rect -96 -48615 -62 -48599
rect 62 -47623 96 -47607
rect 62 -48615 96 -48599
rect -50 -48683 -34 -48649
rect 34 -48683 50 -48649
rect -50 -48791 -34 -48757
rect 34 -48791 50 -48757
rect -96 -48841 -62 -48825
rect -96 -49833 -62 -49817
rect 62 -48841 96 -48825
rect 62 -49833 96 -49817
rect -50 -49901 -34 -49867
rect 34 -49901 50 -49867
rect -50 -50009 -34 -49975
rect 34 -50009 50 -49975
rect -96 -50059 -62 -50043
rect -96 -51051 -62 -51035
rect 62 -50059 96 -50043
rect 62 -51051 96 -51035
rect -50 -51119 -34 -51085
rect 34 -51119 50 -51085
rect -50 -51227 -34 -51193
rect 34 -51227 50 -51193
rect -96 -51277 -62 -51261
rect -96 -52269 -62 -52253
rect 62 -51277 96 -51261
rect 62 -52269 96 -52253
rect -50 -52337 -34 -52303
rect 34 -52337 50 -52303
rect -50 -52445 -34 -52411
rect 34 -52445 50 -52411
rect -96 -52495 -62 -52479
rect -96 -53487 -62 -53471
rect 62 -52495 96 -52479
rect 62 -53487 96 -53471
rect -50 -53555 -34 -53521
rect 34 -53555 50 -53521
rect -50 -53663 -34 -53629
rect 34 -53663 50 -53629
rect -96 -53713 -62 -53697
rect -96 -54705 -62 -54689
rect 62 -53713 96 -53697
rect 62 -54705 96 -54689
rect -50 -54773 -34 -54739
rect 34 -54773 50 -54739
rect -50 -54881 -34 -54847
rect 34 -54881 50 -54847
rect -96 -54931 -62 -54915
rect -96 -55923 -62 -55907
rect 62 -54931 96 -54915
rect 62 -55923 96 -55907
rect -50 -55991 -34 -55957
rect 34 -55991 50 -55957
rect -50 -56099 -34 -56065
rect 34 -56099 50 -56065
rect -96 -56149 -62 -56133
rect -96 -57141 -62 -57125
rect 62 -56149 96 -56133
rect 62 -57141 96 -57125
rect -50 -57209 -34 -57175
rect 34 -57209 50 -57175
rect -50 -57317 -34 -57283
rect 34 -57317 50 -57283
rect -96 -57367 -62 -57351
rect -96 -58359 -62 -58343
rect 62 -57367 96 -57351
rect 62 -58359 96 -58343
rect -50 -58427 -34 -58393
rect 34 -58427 50 -58393
rect -50 -58535 -34 -58501
rect 34 -58535 50 -58501
rect -96 -58585 -62 -58569
rect -96 -59577 -62 -59561
rect 62 -58585 96 -58569
rect 62 -59577 96 -59561
rect -50 -59645 -34 -59611
rect 34 -59645 50 -59611
rect -50 -59753 -34 -59719
rect 34 -59753 50 -59719
rect -96 -59803 -62 -59787
rect -96 -60795 -62 -60779
rect 62 -59803 96 -59787
rect 62 -60795 96 -60779
rect -50 -60863 -34 -60829
rect 34 -60863 50 -60829
rect -50 -60971 -34 -60937
rect 34 -60971 50 -60937
rect -96 -61021 -62 -61005
rect -96 -62013 -62 -61997
rect 62 -61021 96 -61005
rect 62 -62013 96 -61997
rect -50 -62081 -34 -62047
rect 34 -62081 50 -62047
rect -50 -62189 -34 -62155
rect 34 -62189 50 -62155
rect -96 -62239 -62 -62223
rect -96 -63231 -62 -63215
rect 62 -62239 96 -62223
rect 62 -63231 96 -63215
rect -50 -63299 -34 -63265
rect 34 -63299 50 -63265
rect -50 -63407 -34 -63373
rect 34 -63407 50 -63373
rect -96 -63457 -62 -63441
rect -96 -64449 -62 -64433
rect 62 -63457 96 -63441
rect 62 -64449 96 -64433
rect -50 -64517 -34 -64483
rect 34 -64517 50 -64483
rect -50 -64625 -34 -64591
rect 34 -64625 50 -64591
rect -96 -64675 -62 -64659
rect -96 -65667 -62 -65651
rect 62 -64675 96 -64659
rect 62 -65667 96 -65651
rect -50 -65735 -34 -65701
rect 34 -65735 50 -65701
rect -50 -65843 -34 -65809
rect 34 -65843 50 -65809
rect -96 -65893 -62 -65877
rect -96 -66885 -62 -66869
rect 62 -65893 96 -65877
rect 62 -66885 96 -66869
rect -50 -66953 -34 -66919
rect 34 -66953 50 -66919
rect -50 -67061 -34 -67027
rect 34 -67061 50 -67027
rect -96 -67111 -62 -67095
rect -96 -68103 -62 -68087
rect 62 -67111 96 -67095
rect 62 -68103 96 -68087
rect -50 -68171 -34 -68137
rect 34 -68171 50 -68137
rect -50 -68279 -34 -68245
rect 34 -68279 50 -68245
rect -96 -68329 -62 -68313
rect -96 -69321 -62 -69305
rect 62 -68329 96 -68313
rect 62 -69321 96 -69305
rect -50 -69389 -34 -69355
rect 34 -69389 50 -69355
rect -50 -69497 -34 -69463
rect 34 -69497 50 -69463
rect -96 -69547 -62 -69531
rect -96 -70539 -62 -70523
rect 62 -69547 96 -69531
rect 62 -70539 96 -70523
rect -50 -70607 -34 -70573
rect 34 -70607 50 -70573
rect -50 -70715 -34 -70681
rect 34 -70715 50 -70681
rect -96 -70765 -62 -70749
rect -96 -71757 -62 -71741
rect 62 -70765 96 -70749
rect 62 -71757 96 -71741
rect -50 -71825 -34 -71791
rect 34 -71825 50 -71791
rect -50 -71933 -34 -71899
rect 34 -71933 50 -71899
rect -96 -71983 -62 -71967
rect -96 -72975 -62 -72959
rect 62 -71983 96 -71967
rect 62 -72975 96 -72959
rect -50 -73043 -34 -73009
rect 34 -73043 50 -73009
rect -50 -73151 -34 -73117
rect 34 -73151 50 -73117
rect -96 -73201 -62 -73185
rect -96 -74193 -62 -74177
rect 62 -73201 96 -73185
rect 62 -74193 96 -74177
rect -50 -74261 -34 -74227
rect 34 -74261 50 -74227
rect -50 -74369 -34 -74335
rect 34 -74369 50 -74335
rect -96 -74419 -62 -74403
rect -96 -75411 -62 -75395
rect 62 -74419 96 -74403
rect 62 -75411 96 -75395
rect -50 -75479 -34 -75445
rect 34 -75479 50 -75445
rect -50 -75587 -34 -75553
rect 34 -75587 50 -75553
rect -96 -75637 -62 -75621
rect -96 -76629 -62 -76613
rect 62 -75637 96 -75621
rect 62 -76629 96 -76613
rect -50 -76697 -34 -76663
rect 34 -76697 50 -76663
rect -50 -76805 -34 -76771
rect 34 -76805 50 -76771
rect -96 -76855 -62 -76839
rect -96 -77847 -62 -77831
rect 62 -76855 96 -76839
rect 62 -77847 96 -77831
rect -50 -77915 -34 -77881
rect 34 -77915 50 -77881
rect -50 -78023 -34 -77989
rect 34 -78023 50 -77989
rect -96 -78073 -62 -78057
rect -96 -79065 -62 -79049
rect 62 -78073 96 -78057
rect 62 -79065 96 -79049
rect -50 -79133 -34 -79099
rect 34 -79133 50 -79099
rect -50 -79241 -34 -79207
rect 34 -79241 50 -79207
rect -96 -79291 -62 -79275
rect -96 -80283 -62 -80267
rect 62 -79291 96 -79275
rect 62 -80283 96 -80267
rect -50 -80351 -34 -80317
rect 34 -80351 50 -80317
rect -50 -80459 -34 -80425
rect 34 -80459 50 -80425
rect -96 -80509 -62 -80493
rect -96 -81501 -62 -81485
rect 62 -80509 96 -80493
rect 62 -81501 96 -81485
rect -50 -81569 -34 -81535
rect 34 -81569 50 -81535
rect -50 -81677 -34 -81643
rect 34 -81677 50 -81643
rect -96 -81727 -62 -81711
rect -96 -82719 -62 -82703
rect 62 -81727 96 -81711
rect 62 -82719 96 -82703
rect -50 -82787 -34 -82753
rect 34 -82787 50 -82753
rect -50 -82895 -34 -82861
rect 34 -82895 50 -82861
rect -96 -82945 -62 -82929
rect -96 -83937 -62 -83921
rect 62 -82945 96 -82929
rect 62 -83937 96 -83921
rect -50 -84005 -34 -83971
rect 34 -84005 50 -83971
rect -50 -84113 -34 -84079
rect 34 -84113 50 -84079
rect -96 -84163 -62 -84147
rect -96 -85155 -62 -85139
rect 62 -84163 96 -84147
rect 62 -85155 96 -85139
rect -50 -85223 -34 -85189
rect 34 -85223 50 -85189
rect -50 -85331 -34 -85297
rect 34 -85331 50 -85297
rect -96 -85381 -62 -85365
rect -96 -86373 -62 -86357
rect 62 -85381 96 -85365
rect 62 -86373 96 -86357
rect -50 -86441 -34 -86407
rect 34 -86441 50 -86407
rect -50 -86549 -34 -86515
rect 34 -86549 50 -86515
rect -96 -86599 -62 -86583
rect -96 -87591 -62 -87575
rect 62 -86599 96 -86583
rect 62 -87591 96 -87575
rect -50 -87659 -34 -87625
rect 34 -87659 50 -87625
rect -50 -87767 -34 -87733
rect 34 -87767 50 -87733
rect -96 -87817 -62 -87801
rect -96 -88809 -62 -88793
rect 62 -87817 96 -87801
rect 62 -88809 96 -88793
rect -50 -88877 -34 -88843
rect 34 -88877 50 -88843
rect -50 -88985 -34 -88951
rect 34 -88985 50 -88951
rect -96 -89035 -62 -89019
rect -96 -90027 -62 -90011
rect 62 -89035 96 -89019
rect 62 -90027 96 -90011
rect -50 -90095 -34 -90061
rect 34 -90095 50 -90061
rect -50 -90203 -34 -90169
rect 34 -90203 50 -90169
rect -96 -90253 -62 -90237
rect -96 -91245 -62 -91229
rect 62 -90253 96 -90237
rect 62 -91245 96 -91229
rect -50 -91313 -34 -91279
rect 34 -91313 50 -91279
rect -50 -91421 -34 -91387
rect 34 -91421 50 -91387
rect -96 -91471 -62 -91455
rect -96 -92463 -62 -92447
rect 62 -91471 96 -91455
rect 62 -92463 96 -92447
rect -50 -92531 -34 -92497
rect 34 -92531 50 -92497
rect -50 -92639 -34 -92605
rect 34 -92639 50 -92605
rect -96 -92689 -62 -92673
rect -96 -93681 -62 -93665
rect 62 -92689 96 -92673
rect 62 -93681 96 -93665
rect -50 -93749 -34 -93715
rect 34 -93749 50 -93715
rect -50 -93857 -34 -93823
rect 34 -93857 50 -93823
rect -96 -93907 -62 -93891
rect -96 -94899 -62 -94883
rect 62 -93907 96 -93891
rect 62 -94899 96 -94883
rect -50 -94967 -34 -94933
rect 34 -94967 50 -94933
rect -50 -95075 -34 -95041
rect 34 -95075 50 -95041
rect -96 -95125 -62 -95109
rect -96 -96117 -62 -96101
rect 62 -95125 96 -95109
rect 62 -96117 96 -96101
rect -50 -96185 -34 -96151
rect 34 -96185 50 -96151
rect -50 -96293 -34 -96259
rect 34 -96293 50 -96259
rect -96 -96343 -62 -96327
rect -96 -97335 -62 -97319
rect 62 -96343 96 -96327
rect 62 -97335 96 -97319
rect -50 -97403 -34 -97369
rect 34 -97403 50 -97369
rect -50 -97511 -34 -97477
rect 34 -97511 50 -97477
rect -96 -97561 -62 -97545
rect -96 -98553 -62 -98537
rect 62 -97561 96 -97545
rect 62 -98553 96 -98537
rect -50 -98621 -34 -98587
rect 34 -98621 50 -98587
rect -50 -98729 -34 -98695
rect 34 -98729 50 -98695
rect -96 -98779 -62 -98763
rect -96 -99771 -62 -99755
rect 62 -98779 96 -98763
rect 62 -99771 96 -99755
rect -50 -99839 -34 -99805
rect 34 -99839 50 -99805
rect -50 -99947 -34 -99913
rect 34 -99947 50 -99913
rect -96 -99997 -62 -99981
rect -96 -100989 -62 -100973
rect 62 -99997 96 -99981
rect 62 -100989 96 -100973
rect -50 -101057 -34 -101023
rect 34 -101057 50 -101023
rect -50 -101165 -34 -101131
rect 34 -101165 50 -101131
rect -96 -101215 -62 -101199
rect -96 -102207 -62 -102191
rect 62 -101215 96 -101199
rect 62 -102207 96 -102191
rect -50 -102275 -34 -102241
rect 34 -102275 50 -102241
rect -50 -102383 -34 -102349
rect 34 -102383 50 -102349
rect -96 -102433 -62 -102417
rect -96 -103425 -62 -103409
rect 62 -102433 96 -102417
rect 62 -103425 96 -103409
rect -50 -103493 -34 -103459
rect 34 -103493 50 -103459
rect -50 -103601 -34 -103567
rect 34 -103601 50 -103567
rect -96 -103651 -62 -103635
rect -96 -104643 -62 -104627
rect 62 -103651 96 -103635
rect 62 -104643 96 -104627
rect -50 -104711 -34 -104677
rect 34 -104711 50 -104677
rect -50 -104819 -34 -104785
rect 34 -104819 50 -104785
rect -96 -104869 -62 -104853
rect -96 -105861 -62 -105845
rect 62 -104869 96 -104853
rect 62 -105861 96 -105845
rect -50 -105929 -34 -105895
rect 34 -105929 50 -105895
rect -50 -106037 -34 -106003
rect 34 -106037 50 -106003
rect -96 -106087 -62 -106071
rect -96 -107079 -62 -107063
rect 62 -106087 96 -106071
rect 62 -107079 96 -107063
rect -50 -107147 -34 -107113
rect 34 -107147 50 -107113
rect -50 -107255 -34 -107221
rect 34 -107255 50 -107221
rect -96 -107305 -62 -107289
rect -96 -108297 -62 -108281
rect 62 -107305 96 -107289
rect 62 -108297 96 -108281
rect -50 -108365 -34 -108331
rect 34 -108365 50 -108331
rect -50 -108473 -34 -108439
rect 34 -108473 50 -108439
rect -96 -108523 -62 -108507
rect -96 -109515 -62 -109499
rect 62 -108523 96 -108507
rect 62 -109515 96 -109499
rect -50 -109583 -34 -109549
rect 34 -109583 50 -109549
rect -50 -109691 -34 -109657
rect 34 -109691 50 -109657
rect -96 -109741 -62 -109725
rect -96 -110733 -62 -110717
rect 62 -109741 96 -109725
rect 62 -110733 96 -110717
rect -50 -110801 -34 -110767
rect 34 -110801 50 -110767
rect -50 -110909 -34 -110875
rect 34 -110909 50 -110875
rect -96 -110959 -62 -110943
rect -96 -111951 -62 -111935
rect 62 -110959 96 -110943
rect 62 -111951 96 -111935
rect -50 -112019 -34 -111985
rect 34 -112019 50 -111985
rect -50 -112127 -34 -112093
rect 34 -112127 50 -112093
rect -96 -112177 -62 -112161
rect -96 -113169 -62 -113153
rect 62 -112177 96 -112161
rect 62 -113169 96 -113153
rect -50 -113237 -34 -113203
rect 34 -113237 50 -113203
rect -50 -113345 -34 -113311
rect 34 -113345 50 -113311
rect -96 -113395 -62 -113379
rect -96 -114387 -62 -114371
rect 62 -113395 96 -113379
rect 62 -114387 96 -114371
rect -50 -114455 -34 -114421
rect 34 -114455 50 -114421
rect -50 -114563 -34 -114529
rect 34 -114563 50 -114529
rect -96 -114613 -62 -114597
rect -96 -115605 -62 -115589
rect 62 -114613 96 -114597
rect 62 -115605 96 -115589
rect -50 -115673 -34 -115639
rect 34 -115673 50 -115639
rect -50 -115781 -34 -115747
rect 34 -115781 50 -115747
rect -96 -115831 -62 -115815
rect -96 -116823 -62 -116807
rect 62 -115831 96 -115815
rect 62 -116823 96 -116807
rect -50 -116891 -34 -116857
rect 34 -116891 50 -116857
rect -50 -116999 -34 -116965
rect 34 -116999 50 -116965
rect -96 -117049 -62 -117033
rect -96 -118041 -62 -118025
rect 62 -117049 96 -117033
rect 62 -118041 96 -118025
rect -50 -118109 -34 -118075
rect 34 -118109 50 -118075
rect -50 -118217 -34 -118183
rect 34 -118217 50 -118183
rect -96 -118267 -62 -118251
rect -96 -119259 -62 -119243
rect 62 -118267 96 -118251
rect 62 -119259 96 -119243
rect -50 -119327 -34 -119293
rect 34 -119327 50 -119293
rect -50 -119435 -34 -119401
rect 34 -119435 50 -119401
rect -96 -119485 -62 -119469
rect -96 -120477 -62 -120461
rect 62 -119485 96 -119469
rect 62 -120477 96 -120461
rect -50 -120545 -34 -120511
rect 34 -120545 50 -120511
rect -50 -120653 -34 -120619
rect 34 -120653 50 -120619
rect -96 -120703 -62 -120687
rect -96 -121695 -62 -121679
rect 62 -120703 96 -120687
rect 62 -121695 96 -121679
rect -50 -121763 -34 -121729
rect 34 -121763 50 -121729
rect -50 -121871 -34 -121837
rect 34 -121871 50 -121837
rect -96 -121921 -62 -121905
rect -96 -122913 -62 -122897
rect 62 -121921 96 -121905
rect 62 -122913 96 -122897
rect -50 -122981 -34 -122947
rect 34 -122981 50 -122947
rect -50 -123089 -34 -123055
rect 34 -123089 50 -123055
rect -96 -123139 -62 -123123
rect -96 -124131 -62 -124115
rect 62 -123139 96 -123123
rect 62 -124131 96 -124115
rect -50 -124199 -34 -124165
rect 34 -124199 50 -124165
rect -50 -124307 -34 -124273
rect 34 -124307 50 -124273
rect -96 -124357 -62 -124341
rect -96 -125349 -62 -125333
rect 62 -124357 96 -124341
rect 62 -125349 96 -125333
rect -50 -125417 -34 -125383
rect 34 -125417 50 -125383
rect -50 -125525 -34 -125491
rect 34 -125525 50 -125491
rect -96 -125575 -62 -125559
rect -96 -126567 -62 -126551
rect 62 -125575 96 -125559
rect 62 -126567 96 -126551
rect -50 -126635 -34 -126601
rect 34 -126635 50 -126601
rect -50 -126743 -34 -126709
rect 34 -126743 50 -126709
rect -96 -126793 -62 -126777
rect -96 -127785 -62 -127769
rect 62 -126793 96 -126777
rect 62 -127785 96 -127769
rect -50 -127853 -34 -127819
rect 34 -127853 50 -127819
rect -50 -127961 -34 -127927
rect 34 -127961 50 -127927
rect -96 -128011 -62 -127995
rect -96 -129003 -62 -128987
rect 62 -128011 96 -127995
rect 62 -129003 96 -128987
rect -50 -129071 -34 -129037
rect 34 -129071 50 -129037
rect -50 -129179 -34 -129145
rect 34 -129179 50 -129145
rect -96 -129229 -62 -129213
rect -96 -130221 -62 -130205
rect 62 -129229 96 -129213
rect 62 -130221 96 -130205
rect -50 -130289 -34 -130255
rect 34 -130289 50 -130255
rect -50 -130397 -34 -130363
rect 34 -130397 50 -130363
rect -96 -130447 -62 -130431
rect -96 -131439 -62 -131423
rect 62 -130447 96 -130431
rect 62 -131439 96 -131423
rect -50 -131507 -34 -131473
rect 34 -131507 50 -131473
rect -50 -131615 -34 -131581
rect 34 -131615 50 -131581
rect -96 -131665 -62 -131649
rect -96 -132657 -62 -132641
rect 62 -131665 96 -131649
rect 62 -132657 96 -132641
rect -50 -132725 -34 -132691
rect 34 -132725 50 -132691
rect -50 -132833 -34 -132799
rect 34 -132833 50 -132799
rect -96 -132883 -62 -132867
rect -96 -133875 -62 -133859
rect 62 -132883 96 -132867
rect 62 -133875 96 -133859
rect -50 -133943 -34 -133909
rect 34 -133943 50 -133909
rect -50 -134051 -34 -134017
rect 34 -134051 50 -134017
rect -96 -134101 -62 -134085
rect -96 -135093 -62 -135077
rect 62 -134101 96 -134085
rect 62 -135093 96 -135077
rect -50 -135161 -34 -135127
rect 34 -135161 50 -135127
rect -50 -135269 -34 -135235
rect 34 -135269 50 -135235
rect -96 -135319 -62 -135303
rect -96 -136311 -62 -136295
rect 62 -135319 96 -135303
rect 62 -136311 96 -136295
rect -50 -136379 -34 -136345
rect 34 -136379 50 -136345
rect -50 -136487 -34 -136453
rect 34 -136487 50 -136453
rect -96 -136537 -62 -136521
rect -96 -137529 -62 -137513
rect 62 -136537 96 -136521
rect 62 -137529 96 -137513
rect -50 -137597 -34 -137563
rect 34 -137597 50 -137563
rect -50 -137705 -34 -137671
rect 34 -137705 50 -137671
rect -96 -137755 -62 -137739
rect -96 -138747 -62 -138731
rect 62 -137755 96 -137739
rect 62 -138747 96 -138731
rect -50 -138815 -34 -138781
rect 34 -138815 50 -138781
rect -50 -138923 -34 -138889
rect 34 -138923 50 -138889
rect -96 -138973 -62 -138957
rect -96 -139965 -62 -139949
rect 62 -138973 96 -138957
rect 62 -139965 96 -139949
rect -50 -140033 -34 -139999
rect 34 -140033 50 -139999
rect -50 -140141 -34 -140107
rect 34 -140141 50 -140107
rect -96 -140191 -62 -140175
rect -96 -141183 -62 -141167
rect 62 -140191 96 -140175
rect 62 -141183 96 -141167
rect -50 -141251 -34 -141217
rect 34 -141251 50 -141217
rect -50 -141359 -34 -141325
rect 34 -141359 50 -141325
rect -96 -141409 -62 -141393
rect -96 -142401 -62 -142385
rect 62 -141409 96 -141393
rect 62 -142401 96 -142385
rect -50 -142469 -34 -142435
rect 34 -142469 50 -142435
rect -50 -142577 -34 -142543
rect 34 -142577 50 -142543
rect -96 -142627 -62 -142611
rect -96 -143619 -62 -143603
rect 62 -142627 96 -142611
rect 62 -143619 96 -143603
rect -50 -143687 -34 -143653
rect 34 -143687 50 -143653
rect -50 -143795 -34 -143761
rect 34 -143795 50 -143761
rect -96 -143845 -62 -143829
rect -96 -144837 -62 -144821
rect 62 -143845 96 -143829
rect 62 -144837 96 -144821
rect -50 -144905 -34 -144871
rect 34 -144905 50 -144871
rect -50 -145013 -34 -144979
rect 34 -145013 50 -144979
rect -96 -145063 -62 -145047
rect -96 -146055 -62 -146039
rect 62 -145063 96 -145047
rect 62 -146055 96 -146039
rect -50 -146123 -34 -146089
rect 34 -146123 50 -146089
rect -50 -146231 -34 -146197
rect 34 -146231 50 -146197
rect -96 -146281 -62 -146265
rect -96 -147273 -62 -147257
rect 62 -146281 96 -146265
rect 62 -147273 96 -147257
rect -50 -147341 -34 -147307
rect 34 -147341 50 -147307
rect -50 -147449 -34 -147415
rect 34 -147449 50 -147415
rect -96 -147499 -62 -147483
rect -96 -148491 -62 -148475
rect 62 -147499 96 -147483
rect 62 -148491 96 -148475
rect -50 -148559 -34 -148525
rect 34 -148559 50 -148525
rect -50 -148667 -34 -148633
rect 34 -148667 50 -148633
rect -96 -148717 -62 -148701
rect -96 -149709 -62 -149693
rect 62 -148717 96 -148701
rect 62 -149709 96 -149693
rect -50 -149777 -34 -149743
rect 34 -149777 50 -149743
rect -50 -149885 -34 -149851
rect 34 -149885 50 -149851
rect -96 -149935 -62 -149919
rect -96 -150927 -62 -150911
rect 62 -149935 96 -149919
rect 62 -150927 96 -150911
rect -50 -150995 -34 -150961
rect 34 -150995 50 -150961
rect -50 -151103 -34 -151069
rect 34 -151103 50 -151069
rect -96 -151153 -62 -151137
rect -96 -152145 -62 -152129
rect 62 -151153 96 -151137
rect 62 -152145 96 -152129
rect -50 -152213 -34 -152179
rect 34 -152213 50 -152179
rect -50 -152321 -34 -152287
rect 34 -152321 50 -152287
rect -96 -152371 -62 -152355
rect -96 -153363 -62 -153347
rect 62 -152371 96 -152355
rect 62 -153363 96 -153347
rect -50 -153431 -34 -153397
rect 34 -153431 50 -153397
rect -50 -153539 -34 -153505
rect 34 -153539 50 -153505
rect -96 -153589 -62 -153573
rect -96 -154581 -62 -154565
rect 62 -153589 96 -153573
rect 62 -154581 96 -154565
rect -50 -154649 -34 -154615
rect 34 -154649 50 -154615
rect -50 -154757 -34 -154723
rect 34 -154757 50 -154723
rect -96 -154807 -62 -154791
rect -96 -155799 -62 -155783
rect 62 -154807 96 -154791
rect 62 -155799 96 -155783
rect -50 -155867 -34 -155833
rect 34 -155867 50 -155833
rect -50 -155975 -34 -155941
rect 34 -155975 50 -155941
rect -96 -156025 -62 -156009
rect -96 -157017 -62 -157001
rect 62 -156025 96 -156009
rect 62 -157017 96 -157001
rect -50 -157085 -34 -157051
rect 34 -157085 50 -157051
rect -50 -157193 -34 -157159
rect 34 -157193 50 -157159
rect -96 -157243 -62 -157227
rect -96 -158235 -62 -158219
rect 62 -157243 96 -157227
rect 62 -158235 96 -158219
rect -50 -158303 -34 -158269
rect 34 -158303 50 -158269
rect -50 -158411 -34 -158377
rect 34 -158411 50 -158377
rect -96 -158461 -62 -158445
rect -96 -159453 -62 -159437
rect 62 -158461 96 -158445
rect 62 -159453 96 -159437
rect -50 -159521 -34 -159487
rect 34 -159521 50 -159487
rect -50 -159629 -34 -159595
rect 34 -159629 50 -159595
rect -96 -159679 -62 -159663
rect -96 -160671 -62 -160655
rect 62 -159679 96 -159663
rect 62 -160671 96 -160655
rect -50 -160739 -34 -160705
rect 34 -160739 50 -160705
rect -50 -160847 -34 -160813
rect 34 -160847 50 -160813
rect -96 -160897 -62 -160881
rect -96 -161889 -62 -161873
rect 62 -160897 96 -160881
rect 62 -161889 96 -161873
rect -50 -161957 -34 -161923
rect 34 -161957 50 -161923
rect -50 -162065 -34 -162031
rect 34 -162065 50 -162031
rect -96 -162115 -62 -162099
rect -96 -163107 -62 -163091
rect 62 -162115 96 -162099
rect 62 -163107 96 -163091
rect -50 -163175 -34 -163141
rect 34 -163175 50 -163141
rect -50 -163283 -34 -163249
rect 34 -163283 50 -163249
rect -96 -163333 -62 -163317
rect -96 -164325 -62 -164309
rect 62 -163333 96 -163317
rect 62 -164325 96 -164309
rect -50 -164393 -34 -164359
rect 34 -164393 50 -164359
rect -50 -164501 -34 -164467
rect 34 -164501 50 -164467
rect -96 -164551 -62 -164535
rect -96 -165543 -62 -165527
rect 62 -164551 96 -164535
rect 62 -165543 96 -165527
rect -50 -165611 -34 -165577
rect 34 -165611 50 -165577
rect -50 -165719 -34 -165685
rect 34 -165719 50 -165685
rect -96 -165769 -62 -165753
rect -96 -166761 -62 -166745
rect 62 -165769 96 -165753
rect 62 -166761 96 -166745
rect -50 -166829 -34 -166795
rect 34 -166829 50 -166795
rect -50 -166937 -34 -166903
rect 34 -166937 50 -166903
rect -96 -166987 -62 -166971
rect -96 -167979 -62 -167963
rect 62 -166987 96 -166971
rect 62 -167979 96 -167963
rect -50 -168047 -34 -168013
rect 34 -168047 50 -168013
rect -50 -168155 -34 -168121
rect 34 -168155 50 -168121
rect -96 -168205 -62 -168189
rect -96 -169197 -62 -169181
rect 62 -168205 96 -168189
rect 62 -169197 96 -169181
rect -50 -169265 -34 -169231
rect 34 -169265 50 -169231
rect -50 -169373 -34 -169339
rect 34 -169373 50 -169339
rect -96 -169423 -62 -169407
rect -96 -170415 -62 -170399
rect 62 -169423 96 -169407
rect 62 -170415 96 -170399
rect -50 -170483 -34 -170449
rect 34 -170483 50 -170449
rect -50 -170591 -34 -170557
rect 34 -170591 50 -170557
rect -96 -170641 -62 -170625
rect -96 -171633 -62 -171617
rect 62 -170641 96 -170625
rect 62 -171633 96 -171617
rect -50 -171701 -34 -171667
rect 34 -171701 50 -171667
rect -50 -171809 -34 -171775
rect 34 -171809 50 -171775
rect -96 -171859 -62 -171843
rect -96 -172851 -62 -172835
rect 62 -171859 96 -171843
rect 62 -172851 96 -172835
rect -50 -172919 -34 -172885
rect 34 -172919 50 -172885
rect -50 -173027 -34 -172993
rect 34 -173027 50 -172993
rect -96 -173077 -62 -173061
rect -96 -174069 -62 -174053
rect 62 -173077 96 -173061
rect 62 -174069 96 -174053
rect -50 -174137 -34 -174103
rect 34 -174137 50 -174103
rect -50 -174245 -34 -174211
rect 34 -174245 50 -174211
rect -96 -174295 -62 -174279
rect -96 -175287 -62 -175271
rect 62 -174295 96 -174279
rect 62 -175287 96 -175271
rect -50 -175355 -34 -175321
rect 34 -175355 50 -175321
rect -50 -175463 -34 -175429
rect 34 -175463 50 -175429
rect -96 -175513 -62 -175497
rect -96 -176505 -62 -176489
rect 62 -175513 96 -175497
rect 62 -176505 96 -176489
rect -50 -176573 -34 -176539
rect 34 -176573 50 -176539
rect -50 -176681 -34 -176647
rect 34 -176681 50 -176647
rect -96 -176731 -62 -176715
rect -96 -177723 -62 -177707
rect 62 -176731 96 -176715
rect 62 -177723 96 -177707
rect -50 -177791 -34 -177757
rect 34 -177791 50 -177757
rect -50 -177899 -34 -177865
rect 34 -177899 50 -177865
rect -96 -177949 -62 -177933
rect -96 -178941 -62 -178925
rect 62 -177949 96 -177933
rect 62 -178941 96 -178925
rect -50 -179009 -34 -178975
rect 34 -179009 50 -178975
rect -50 -179117 -34 -179083
rect 34 -179117 50 -179083
rect -96 -179167 -62 -179151
rect -96 -180159 -62 -180143
rect 62 -179167 96 -179151
rect 62 -180159 96 -180143
rect -50 -180227 -34 -180193
rect 34 -180227 50 -180193
rect -50 -180335 -34 -180301
rect 34 -180335 50 -180301
rect -96 -180385 -62 -180369
rect -96 -181377 -62 -181361
rect 62 -180385 96 -180369
rect 62 -181377 96 -181361
rect -50 -181445 -34 -181411
rect 34 -181445 50 -181411
rect -50 -181553 -34 -181519
rect 34 -181553 50 -181519
rect -96 -181603 -62 -181587
rect -96 -182595 -62 -182579
rect 62 -181603 96 -181587
rect 62 -182595 96 -182579
rect -50 -182663 -34 -182629
rect 34 -182663 50 -182629
rect -50 -182771 -34 -182737
rect 34 -182771 50 -182737
rect -96 -182821 -62 -182805
rect -96 -183813 -62 -183797
rect 62 -182821 96 -182805
rect 62 -183813 96 -183797
rect -50 -183881 -34 -183847
rect 34 -183881 50 -183847
rect -50 -183989 -34 -183955
rect 34 -183989 50 -183955
rect -96 -184039 -62 -184023
rect -96 -185031 -62 -185015
rect 62 -184039 96 -184023
rect 62 -185031 96 -185015
rect -50 -185099 -34 -185065
rect 34 -185099 50 -185065
rect -50 -185207 -34 -185173
rect 34 -185207 50 -185173
rect -96 -185257 -62 -185241
rect -96 -186249 -62 -186233
rect 62 -185257 96 -185241
rect 62 -186249 96 -186233
rect -50 -186317 -34 -186283
rect 34 -186317 50 -186283
rect -50 -186425 -34 -186391
rect 34 -186425 50 -186391
rect -96 -186475 -62 -186459
rect -96 -187467 -62 -187451
rect 62 -186475 96 -186459
rect 62 -187467 96 -187451
rect -50 -187535 -34 -187501
rect 34 -187535 50 -187501
rect -50 -187643 -34 -187609
rect 34 -187643 50 -187609
rect -96 -187693 -62 -187677
rect -96 -188685 -62 -188669
rect 62 -187693 96 -187677
rect 62 -188685 96 -188669
rect -50 -188753 -34 -188719
rect 34 -188753 50 -188719
rect -50 -188861 -34 -188827
rect 34 -188861 50 -188827
rect -96 -188911 -62 -188895
rect -96 -189903 -62 -189887
rect 62 -188911 96 -188895
rect 62 -189903 96 -189887
rect -50 -189971 -34 -189937
rect 34 -189971 50 -189937
rect -50 -190079 -34 -190045
rect 34 -190079 50 -190045
rect -96 -190129 -62 -190113
rect -96 -191121 -62 -191105
rect 62 -190129 96 -190113
rect 62 -191121 96 -191105
rect -50 -191189 -34 -191155
rect 34 -191189 50 -191155
rect -50 -191297 -34 -191263
rect 34 -191297 50 -191263
rect -96 -191347 -62 -191331
rect -96 -192339 -62 -192323
rect 62 -191347 96 -191331
rect 62 -192339 96 -192323
rect -50 -192407 -34 -192373
rect 34 -192407 50 -192373
rect -50 -192515 -34 -192481
rect 34 -192515 50 -192481
rect -96 -192565 -62 -192549
rect -96 -193557 -62 -193541
rect 62 -192565 96 -192549
rect 62 -193557 96 -193541
rect -50 -193625 -34 -193591
rect 34 -193625 50 -193591
rect -50 -193733 -34 -193699
rect 34 -193733 50 -193699
rect -96 -193783 -62 -193767
rect -96 -194775 -62 -194759
rect 62 -193783 96 -193767
rect 62 -194775 96 -194759
rect -50 -194843 -34 -194809
rect 34 -194843 50 -194809
rect -50 -194951 -34 -194917
rect 34 -194951 50 -194917
rect -96 -195001 -62 -194985
rect -96 -195993 -62 -195977
rect 62 -195001 96 -194985
rect 62 -195993 96 -195977
rect -50 -196061 -34 -196027
rect 34 -196061 50 -196027
rect -50 -196169 -34 -196135
rect 34 -196169 50 -196135
rect -96 -196219 -62 -196203
rect -96 -197211 -62 -197195
rect 62 -196219 96 -196203
rect 62 -197211 96 -197195
rect -50 -197279 -34 -197245
rect 34 -197279 50 -197245
rect -50 -197387 -34 -197353
rect 34 -197387 50 -197353
rect -96 -197437 -62 -197421
rect -96 -198429 -62 -198413
rect 62 -197437 96 -197421
rect 62 -198429 96 -198413
rect -50 -198497 -34 -198463
rect 34 -198497 50 -198463
rect -50 -198605 -34 -198571
rect 34 -198605 50 -198571
rect -96 -198655 -62 -198639
rect -96 -199647 -62 -199631
rect 62 -198655 96 -198639
rect 62 -199647 96 -199631
rect -50 -199715 -34 -199681
rect 34 -199715 50 -199681
rect -50 -199823 -34 -199789
rect 34 -199823 50 -199789
rect -96 -199873 -62 -199857
rect -96 -200865 -62 -200849
rect 62 -199873 96 -199857
rect 62 -200865 96 -200849
rect -50 -200933 -34 -200899
rect 34 -200933 50 -200899
rect -50 -201041 -34 -201007
rect 34 -201041 50 -201007
rect -96 -201091 -62 -201075
rect -96 -202083 -62 -202067
rect 62 -201091 96 -201075
rect 62 -202083 96 -202067
rect -50 -202151 -34 -202117
rect 34 -202151 50 -202117
rect -50 -202259 -34 -202225
rect 34 -202259 50 -202225
rect -96 -202309 -62 -202293
rect -96 -203301 -62 -203285
rect 62 -202309 96 -202293
rect 62 -203301 96 -203285
rect -50 -203369 -34 -203335
rect 34 -203369 50 -203335
rect -50 -203477 -34 -203443
rect 34 -203477 50 -203443
rect -96 -203527 -62 -203511
rect -96 -204519 -62 -204503
rect 62 -203527 96 -203511
rect 62 -204519 96 -204503
rect -50 -204587 -34 -204553
rect 34 -204587 50 -204553
rect -50 -204695 -34 -204661
rect 34 -204695 50 -204661
rect -96 -204745 -62 -204729
rect -96 -205737 -62 -205721
rect 62 -204745 96 -204729
rect 62 -205737 96 -205721
rect -50 -205805 -34 -205771
rect 34 -205805 50 -205771
rect -50 -205913 -34 -205879
rect 34 -205913 50 -205879
rect -96 -205963 -62 -205947
rect -96 -206955 -62 -206939
rect 62 -205963 96 -205947
rect 62 -206955 96 -206939
rect -50 -207023 -34 -206989
rect 34 -207023 50 -206989
rect -50 -207131 -34 -207097
rect 34 -207131 50 -207097
rect -96 -207181 -62 -207165
rect -96 -208173 -62 -208157
rect 62 -207181 96 -207165
rect 62 -208173 96 -208157
rect -50 -208241 -34 -208207
rect 34 -208241 50 -208207
rect -50 -208349 -34 -208315
rect 34 -208349 50 -208315
rect -96 -208399 -62 -208383
rect -96 -209391 -62 -209375
rect 62 -208399 96 -208383
rect 62 -209391 96 -209375
rect -50 -209459 -34 -209425
rect 34 -209459 50 -209425
rect -50 -209567 -34 -209533
rect 34 -209567 50 -209533
rect -96 -209617 -62 -209601
rect -96 -210609 -62 -210593
rect 62 -209617 96 -209601
rect 62 -210609 96 -210593
rect -50 -210677 -34 -210643
rect 34 -210677 50 -210643
rect -50 -210785 -34 -210751
rect 34 -210785 50 -210751
rect -96 -210835 -62 -210819
rect -96 -211827 -62 -211811
rect 62 -210835 96 -210819
rect 62 -211827 96 -211811
rect -50 -211895 -34 -211861
rect 34 -211895 50 -211861
rect -50 -212003 -34 -211969
rect 34 -212003 50 -211969
rect -96 -212053 -62 -212037
rect -96 -213045 -62 -213029
rect 62 -212053 96 -212037
rect 62 -213045 96 -213029
rect -50 -213113 -34 -213079
rect 34 -213113 50 -213079
rect -50 -213221 -34 -213187
rect 34 -213221 50 -213187
rect -96 -213271 -62 -213255
rect -96 -214263 -62 -214247
rect 62 -213271 96 -213255
rect 62 -214263 96 -214247
rect -50 -214331 -34 -214297
rect 34 -214331 50 -214297
rect -50 -214439 -34 -214405
rect 34 -214439 50 -214405
rect -96 -214489 -62 -214473
rect -96 -215481 -62 -215465
rect 62 -214489 96 -214473
rect 62 -215481 96 -215465
rect -50 -215549 -34 -215515
rect 34 -215549 50 -215515
rect -50 -215657 -34 -215623
rect 34 -215657 50 -215623
rect -96 -215707 -62 -215691
rect -96 -216699 -62 -216683
rect 62 -215707 96 -215691
rect 62 -216699 96 -216683
rect -50 -216767 -34 -216733
rect 34 -216767 50 -216733
rect -50 -216875 -34 -216841
rect 34 -216875 50 -216841
rect -96 -216925 -62 -216909
rect -96 -217917 -62 -217901
rect 62 -216925 96 -216909
rect 62 -217917 96 -217901
rect -50 -217985 -34 -217951
rect 34 -217985 50 -217951
rect -50 -218093 -34 -218059
rect 34 -218093 50 -218059
rect -96 -218143 -62 -218127
rect -96 -219135 -62 -219119
rect 62 -218143 96 -218127
rect 62 -219135 96 -219119
rect -50 -219203 -34 -219169
rect 34 -219203 50 -219169
rect -50 -219311 -34 -219277
rect 34 -219311 50 -219277
rect -96 -219361 -62 -219345
rect -96 -220353 -62 -220337
rect 62 -219361 96 -219345
rect 62 -220353 96 -220337
rect -50 -220421 -34 -220387
rect 34 -220421 50 -220387
rect -50 -220529 -34 -220495
rect 34 -220529 50 -220495
rect -96 -220579 -62 -220563
rect -96 -221571 -62 -221555
rect 62 -220579 96 -220563
rect 62 -221571 96 -221555
rect -50 -221639 -34 -221605
rect 34 -221639 50 -221605
rect -50 -221747 -34 -221713
rect 34 -221747 50 -221713
rect -96 -221797 -62 -221781
rect -96 -222789 -62 -222773
rect 62 -221797 96 -221781
rect 62 -222789 96 -222773
rect -50 -222857 -34 -222823
rect 34 -222857 50 -222823
rect -50 -222965 -34 -222931
rect 34 -222965 50 -222931
rect -96 -223015 -62 -222999
rect -96 -224007 -62 -223991
rect 62 -223015 96 -222999
rect 62 -224007 96 -223991
rect -50 -224075 -34 -224041
rect 34 -224075 50 -224041
rect -50 -224183 -34 -224149
rect 34 -224183 50 -224149
rect -96 -224233 -62 -224217
rect -96 -225225 -62 -225209
rect 62 -224233 96 -224217
rect 62 -225225 96 -225209
rect -50 -225293 -34 -225259
rect 34 -225293 50 -225259
rect -50 -225401 -34 -225367
rect 34 -225401 50 -225367
rect -96 -225451 -62 -225435
rect -96 -226443 -62 -226427
rect 62 -225451 96 -225435
rect 62 -226443 96 -226427
rect -50 -226511 -34 -226477
rect 34 -226511 50 -226477
rect -50 -226619 -34 -226585
rect 34 -226619 50 -226585
rect -96 -226669 -62 -226653
rect -96 -227661 -62 -227645
rect 62 -226669 96 -226653
rect 62 -227661 96 -227645
rect -50 -227729 -34 -227695
rect 34 -227729 50 -227695
rect -50 -227837 -34 -227803
rect 34 -227837 50 -227803
rect -96 -227887 -62 -227871
rect -96 -228879 -62 -228863
rect 62 -227887 96 -227871
rect 62 -228879 96 -228863
rect -50 -228947 -34 -228913
rect 34 -228947 50 -228913
rect -50 -229055 -34 -229021
rect 34 -229055 50 -229021
rect -96 -229105 -62 -229089
rect -96 -230097 -62 -230081
rect 62 -229105 96 -229089
rect 62 -230097 96 -230081
rect -50 -230165 -34 -230131
rect 34 -230165 50 -230131
rect -50 -230273 -34 -230239
rect 34 -230273 50 -230239
rect -96 -230323 -62 -230307
rect -96 -231315 -62 -231299
rect 62 -230323 96 -230307
rect 62 -231315 96 -231299
rect -50 -231383 -34 -231349
rect 34 -231383 50 -231349
rect -50 -231491 -34 -231457
rect 34 -231491 50 -231457
rect -96 -231541 -62 -231525
rect -96 -232533 -62 -232517
rect 62 -231541 96 -231525
rect 62 -232533 96 -232517
rect -50 -232601 -34 -232567
rect 34 -232601 50 -232567
rect -50 -232709 -34 -232675
rect 34 -232709 50 -232675
rect -96 -232759 -62 -232743
rect -96 -233751 -62 -233735
rect 62 -232759 96 -232743
rect 62 -233751 96 -233735
rect -50 -233819 -34 -233785
rect 34 -233819 50 -233785
rect -50 -233927 -34 -233893
rect 34 -233927 50 -233893
rect -96 -233977 -62 -233961
rect -96 -234969 -62 -234953
rect 62 -233977 96 -233961
rect 62 -234969 96 -234953
rect -50 -235037 -34 -235003
rect 34 -235037 50 -235003
rect -50 -235145 -34 -235111
rect 34 -235145 50 -235111
rect -96 -235195 -62 -235179
rect -96 -236187 -62 -236171
rect 62 -235195 96 -235179
rect 62 -236187 96 -236171
rect -50 -236255 -34 -236221
rect 34 -236255 50 -236221
rect -50 -236363 -34 -236329
rect 34 -236363 50 -236329
rect -96 -236413 -62 -236397
rect -96 -237405 -62 -237389
rect 62 -236413 96 -236397
rect 62 -237405 96 -237389
rect -50 -237473 -34 -237439
rect 34 -237473 50 -237439
rect -50 -237581 -34 -237547
rect 34 -237581 50 -237547
rect -96 -237631 -62 -237615
rect -96 -238623 -62 -238607
rect 62 -237631 96 -237615
rect 62 -238623 96 -238607
rect -50 -238691 -34 -238657
rect 34 -238691 50 -238657
rect -50 -238799 -34 -238765
rect 34 -238799 50 -238765
rect -96 -238849 -62 -238833
rect -96 -239841 -62 -239825
rect 62 -238849 96 -238833
rect 62 -239841 96 -239825
rect -50 -239909 -34 -239875
rect 34 -239909 50 -239875
rect -50 -240017 -34 -239983
rect 34 -240017 50 -239983
rect -96 -240067 -62 -240051
rect -96 -241059 -62 -241043
rect 62 -240067 96 -240051
rect 62 -241059 96 -241043
rect -50 -241127 -34 -241093
rect 34 -241127 50 -241093
rect -50 -241235 -34 -241201
rect 34 -241235 50 -241201
rect -96 -241285 -62 -241269
rect -96 -242277 -62 -242261
rect 62 -241285 96 -241269
rect 62 -242277 96 -242261
rect -50 -242345 -34 -242311
rect 34 -242345 50 -242311
rect -50 -242453 -34 -242419
rect 34 -242453 50 -242419
rect -96 -242503 -62 -242487
rect -96 -243495 -62 -243479
rect 62 -242503 96 -242487
rect 62 -243495 96 -243479
rect -50 -243563 -34 -243529
rect 34 -243563 50 -243529
rect -50 -243671 -34 -243637
rect 34 -243671 50 -243637
rect -96 -243721 -62 -243705
rect -96 -244713 -62 -244697
rect 62 -243721 96 -243705
rect 62 -244713 96 -244697
rect -50 -244781 -34 -244747
rect 34 -244781 50 -244747
rect -50 -244889 -34 -244855
rect 34 -244889 50 -244855
rect -96 -244939 -62 -244923
rect -96 -245931 -62 -245915
rect 62 -244939 96 -244923
rect 62 -245931 96 -245915
rect -50 -245999 -34 -245965
rect 34 -245999 50 -245965
rect -50 -246107 -34 -246073
rect 34 -246107 50 -246073
rect -96 -246157 -62 -246141
rect -96 -247149 -62 -247133
rect 62 -246157 96 -246141
rect 62 -247149 96 -247133
rect -50 -247217 -34 -247183
rect 34 -247217 50 -247183
rect -50 -247325 -34 -247291
rect 34 -247325 50 -247291
rect -96 -247375 -62 -247359
rect -96 -248367 -62 -248351
rect 62 -247375 96 -247359
rect 62 -248367 96 -248351
rect -50 -248435 -34 -248401
rect 34 -248435 50 -248401
rect -50 -248543 -34 -248509
rect 34 -248543 50 -248509
rect -96 -248593 -62 -248577
rect -96 -249585 -62 -249569
rect 62 -248593 96 -248577
rect 62 -249585 96 -249569
rect -50 -249653 -34 -249619
rect 34 -249653 50 -249619
rect -50 -249761 -34 -249727
rect 34 -249761 50 -249727
rect -96 -249811 -62 -249795
rect -96 -250803 -62 -250787
rect 62 -249811 96 -249795
rect 62 -250803 96 -250787
rect -50 -250871 -34 -250837
rect 34 -250871 50 -250837
rect -50 -250979 -34 -250945
rect 34 -250979 50 -250945
rect -96 -251029 -62 -251013
rect -96 -252021 -62 -252005
rect 62 -251029 96 -251013
rect 62 -252021 96 -252005
rect -50 -252089 -34 -252055
rect 34 -252089 50 -252055
rect -50 -252197 -34 -252163
rect 34 -252197 50 -252163
rect -96 -252247 -62 -252231
rect -96 -253239 -62 -253223
rect 62 -252247 96 -252231
rect 62 -253239 96 -253223
rect -50 -253307 -34 -253273
rect 34 -253307 50 -253273
rect -50 -253415 -34 -253381
rect 34 -253415 50 -253381
rect -96 -253465 -62 -253449
rect -96 -254457 -62 -254441
rect 62 -253465 96 -253449
rect 62 -254457 96 -254441
rect -50 -254525 -34 -254491
rect 34 -254525 50 -254491
rect -50 -254633 -34 -254599
rect 34 -254633 50 -254599
rect -96 -254683 -62 -254667
rect -96 -255675 -62 -255659
rect 62 -254683 96 -254667
rect 62 -255675 96 -255659
rect -50 -255743 -34 -255709
rect 34 -255743 50 -255709
rect -50 -255851 -34 -255817
rect 34 -255851 50 -255817
rect -96 -255901 -62 -255885
rect -96 -256893 -62 -256877
rect 62 -255901 96 -255885
rect 62 -256893 96 -256877
rect -50 -256961 -34 -256927
rect 34 -256961 50 -256927
rect -50 -257069 -34 -257035
rect 34 -257069 50 -257035
rect -96 -257119 -62 -257103
rect -96 -258111 -62 -258095
rect 62 -257119 96 -257103
rect 62 -258111 96 -258095
rect -50 -258179 -34 -258145
rect 34 -258179 50 -258145
rect -50 -258287 -34 -258253
rect 34 -258287 50 -258253
rect -96 -258337 -62 -258321
rect -96 -259329 -62 -259313
rect 62 -258337 96 -258321
rect 62 -259329 96 -259313
rect -50 -259397 -34 -259363
rect 34 -259397 50 -259363
rect -50 -259505 -34 -259471
rect 34 -259505 50 -259471
rect -96 -259555 -62 -259539
rect -96 -260547 -62 -260531
rect 62 -259555 96 -259539
rect 62 -260547 96 -260531
rect -50 -260615 -34 -260581
rect 34 -260615 50 -260581
rect -50 -260723 -34 -260689
rect 34 -260723 50 -260689
rect -96 -260773 -62 -260757
rect -96 -261765 -62 -261749
rect 62 -260773 96 -260757
rect 62 -261765 96 -261749
rect -50 -261833 -34 -261799
rect 34 -261833 50 -261799
rect -50 -261941 -34 -261907
rect 34 -261941 50 -261907
rect -96 -261991 -62 -261975
rect -96 -262983 -62 -262967
rect 62 -261991 96 -261975
rect 62 -262983 96 -262967
rect -50 -263051 -34 -263017
rect 34 -263051 50 -263017
rect -50 -263159 -34 -263125
rect 34 -263159 50 -263125
rect -96 -263209 -62 -263193
rect -96 -264201 -62 -264185
rect 62 -263209 96 -263193
rect 62 -264201 96 -264185
rect -50 -264269 -34 -264235
rect 34 -264269 50 -264235
rect -50 -264377 -34 -264343
rect 34 -264377 50 -264343
rect -96 -264427 -62 -264411
rect -96 -265419 -62 -265403
rect 62 -264427 96 -264411
rect 62 -265419 96 -265403
rect -50 -265487 -34 -265453
rect 34 -265487 50 -265453
rect -50 -265595 -34 -265561
rect 34 -265595 50 -265561
rect -96 -265645 -62 -265629
rect -96 -266637 -62 -266621
rect 62 -265645 96 -265629
rect 62 -266637 96 -266621
rect -50 -266705 -34 -266671
rect 34 -266705 50 -266671
rect -50 -266813 -34 -266779
rect 34 -266813 50 -266779
rect -96 -266863 -62 -266847
rect -96 -267855 -62 -267839
rect 62 -266863 96 -266847
rect 62 -267855 96 -267839
rect -50 -267923 -34 -267889
rect 34 -267923 50 -267889
rect -50 -268031 -34 -267997
rect 34 -268031 50 -267997
rect -96 -268081 -62 -268065
rect -96 -269073 -62 -269057
rect 62 -268081 96 -268065
rect 62 -269073 96 -269057
rect -50 -269141 -34 -269107
rect 34 -269141 50 -269107
rect -50 -269249 -34 -269215
rect 34 -269249 50 -269215
rect -96 -269299 -62 -269283
rect -96 -270291 -62 -270275
rect 62 -269299 96 -269283
rect 62 -270291 96 -270275
rect -50 -270359 -34 -270325
rect 34 -270359 50 -270325
rect -50 -270467 -34 -270433
rect 34 -270467 50 -270433
rect -96 -270517 -62 -270501
rect -96 -271509 -62 -271493
rect 62 -270517 96 -270501
rect 62 -271509 96 -271493
rect -50 -271577 -34 -271543
rect 34 -271577 50 -271543
rect -50 -271685 -34 -271651
rect 34 -271685 50 -271651
rect -96 -271735 -62 -271719
rect -96 -272727 -62 -272711
rect 62 -271735 96 -271719
rect 62 -272727 96 -272711
rect -50 -272795 -34 -272761
rect 34 -272795 50 -272761
rect -50 -272903 -34 -272869
rect 34 -272903 50 -272869
rect -96 -272953 -62 -272937
rect -96 -273945 -62 -273929
rect 62 -272953 96 -272937
rect 62 -273945 96 -273929
rect -50 -274013 -34 -273979
rect 34 -274013 50 -273979
rect -50 -274121 -34 -274087
rect 34 -274121 50 -274087
rect -96 -274171 -62 -274155
rect -96 -275163 -62 -275147
rect 62 -274171 96 -274155
rect 62 -275163 96 -275147
rect -50 -275231 -34 -275197
rect 34 -275231 50 -275197
rect -50 -275339 -34 -275305
rect 34 -275339 50 -275305
rect -96 -275389 -62 -275373
rect -96 -276381 -62 -276365
rect 62 -275389 96 -275373
rect 62 -276381 96 -276365
rect -50 -276449 -34 -276415
rect 34 -276449 50 -276415
rect -50 -276557 -34 -276523
rect 34 -276557 50 -276523
rect -96 -276607 -62 -276591
rect -96 -277599 -62 -277583
rect 62 -276607 96 -276591
rect 62 -277599 96 -277583
rect -50 -277667 -34 -277633
rect 34 -277667 50 -277633
rect -50 -277775 -34 -277741
rect 34 -277775 50 -277741
rect -96 -277825 -62 -277809
rect -96 -278817 -62 -278801
rect 62 -277825 96 -277809
rect 62 -278817 96 -278801
rect -50 -278885 -34 -278851
rect 34 -278885 50 -278851
rect -50 -278993 -34 -278959
rect 34 -278993 50 -278959
rect -96 -279043 -62 -279027
rect -96 -280035 -62 -280019
rect 62 -279043 96 -279027
rect 62 -280035 96 -280019
rect -50 -280103 -34 -280069
rect 34 -280103 50 -280069
rect -50 -280211 -34 -280177
rect 34 -280211 50 -280177
rect -96 -280261 -62 -280245
rect -96 -281253 -62 -281237
rect 62 -280261 96 -280245
rect 62 -281253 96 -281237
rect -50 -281321 -34 -281287
rect 34 -281321 50 -281287
rect -50 -281429 -34 -281395
rect 34 -281429 50 -281395
rect -96 -281479 -62 -281463
rect -96 -282471 -62 -282455
rect 62 -281479 96 -281463
rect 62 -282471 96 -282455
rect -50 -282539 -34 -282505
rect 34 -282539 50 -282505
rect -50 -282647 -34 -282613
rect 34 -282647 50 -282613
rect -96 -282697 -62 -282681
rect -96 -283689 -62 -283673
rect 62 -282697 96 -282681
rect 62 -283689 96 -283673
rect -50 -283757 -34 -283723
rect 34 -283757 50 -283723
rect -50 -283865 -34 -283831
rect 34 -283865 50 -283831
rect -96 -283915 -62 -283899
rect -96 -284907 -62 -284891
rect 62 -283915 96 -283899
rect 62 -284907 96 -284891
rect -50 -284975 -34 -284941
rect 34 -284975 50 -284941
rect -50 -285083 -34 -285049
rect 34 -285083 50 -285049
rect -96 -285133 -62 -285117
rect -96 -286125 -62 -286109
rect 62 -285133 96 -285117
rect 62 -286125 96 -286109
rect -50 -286193 -34 -286159
rect 34 -286193 50 -286159
rect -50 -286301 -34 -286267
rect 34 -286301 50 -286267
rect -96 -286351 -62 -286335
rect -96 -287343 -62 -287327
rect 62 -286351 96 -286335
rect 62 -287343 96 -287327
rect -50 -287411 -34 -287377
rect 34 -287411 50 -287377
rect -50 -287519 -34 -287485
rect 34 -287519 50 -287485
rect -96 -287569 -62 -287553
rect -96 -288561 -62 -288545
rect 62 -287569 96 -287553
rect 62 -288561 96 -288545
rect -50 -288629 -34 -288595
rect 34 -288629 50 -288595
rect -50 -288737 -34 -288703
rect 34 -288737 50 -288703
rect -96 -288787 -62 -288771
rect -96 -289779 -62 -289763
rect 62 -288787 96 -288771
rect 62 -289779 96 -289763
rect -50 -289847 -34 -289813
rect 34 -289847 50 -289813
rect -50 -289955 -34 -289921
rect 34 -289955 50 -289921
rect -96 -290005 -62 -289989
rect -96 -290997 -62 -290981
rect 62 -290005 96 -289989
rect 62 -290997 96 -290981
rect -50 -291065 -34 -291031
rect 34 -291065 50 -291031
rect -50 -291173 -34 -291139
rect 34 -291173 50 -291139
rect -96 -291223 -62 -291207
rect -96 -292215 -62 -292199
rect 62 -291223 96 -291207
rect 62 -292215 96 -292199
rect -50 -292283 -34 -292249
rect 34 -292283 50 -292249
rect -50 -292391 -34 -292357
rect 34 -292391 50 -292357
rect -96 -292441 -62 -292425
rect -96 -293433 -62 -293417
rect 62 -292441 96 -292425
rect 62 -293433 96 -293417
rect -50 -293501 -34 -293467
rect 34 -293501 50 -293467
rect -50 -293609 -34 -293575
rect 34 -293609 50 -293575
rect -96 -293659 -62 -293643
rect -96 -294651 -62 -294635
rect 62 -293659 96 -293643
rect 62 -294651 96 -294635
rect -50 -294719 -34 -294685
rect 34 -294719 50 -294685
rect -50 -294827 -34 -294793
rect 34 -294827 50 -294793
rect -96 -294877 -62 -294861
rect -96 -295869 -62 -295853
rect 62 -294877 96 -294861
rect 62 -295869 96 -295853
rect -50 -295937 -34 -295903
rect 34 -295937 50 -295903
rect -50 -296045 -34 -296011
rect 34 -296045 50 -296011
rect -96 -296095 -62 -296079
rect -96 -297087 -62 -297071
rect 62 -296095 96 -296079
rect 62 -297087 96 -297071
rect -50 -297155 -34 -297121
rect 34 -297155 50 -297121
rect -50 -297263 -34 -297229
rect 34 -297263 50 -297229
rect -96 -297313 -62 -297297
rect -96 -298305 -62 -298289
rect 62 -297313 96 -297297
rect 62 -298305 96 -298289
rect -50 -298373 -34 -298339
rect 34 -298373 50 -298339
rect -50 -298481 -34 -298447
rect 34 -298481 50 -298447
rect -96 -298531 -62 -298515
rect -96 -299523 -62 -299507
rect 62 -298531 96 -298515
rect 62 -299523 96 -299507
rect -50 -299591 -34 -299557
rect 34 -299591 50 -299557
rect -50 -299699 -34 -299665
rect 34 -299699 50 -299665
rect -96 -299749 -62 -299733
rect -96 -300741 -62 -300725
rect 62 -299749 96 -299733
rect 62 -300741 96 -300725
rect -50 -300809 -34 -300775
rect 34 -300809 50 -300775
rect -50 -300917 -34 -300883
rect 34 -300917 50 -300883
rect -96 -300967 -62 -300951
rect -96 -301959 -62 -301943
rect 62 -300967 96 -300951
rect 62 -301959 96 -301943
rect -50 -302027 -34 -301993
rect 34 -302027 50 -301993
rect -50 -302135 -34 -302101
rect 34 -302135 50 -302101
rect -96 -302185 -62 -302169
rect -96 -303177 -62 -303161
rect 62 -302185 96 -302169
rect 62 -303177 96 -303161
rect -50 -303245 -34 -303211
rect 34 -303245 50 -303211
rect -50 -303353 -34 -303319
rect 34 -303353 50 -303319
rect -96 -303403 -62 -303387
rect -96 -304395 -62 -304379
rect 62 -303403 96 -303387
rect 62 -304395 96 -304379
rect -50 -304463 -34 -304429
rect 34 -304463 50 -304429
rect -50 -304571 -34 -304537
rect 34 -304571 50 -304537
rect -96 -304621 -62 -304605
rect -96 -305613 -62 -305597
rect 62 -304621 96 -304605
rect 62 -305613 96 -305597
rect -50 -305681 -34 -305647
rect 34 -305681 50 -305647
rect -50 -305789 -34 -305755
rect 34 -305789 50 -305755
rect -96 -305839 -62 -305823
rect -96 -306831 -62 -306815
rect 62 -305839 96 -305823
rect 62 -306831 96 -306815
rect -50 -306899 -34 -306865
rect 34 -306899 50 -306865
rect -50 -307007 -34 -306973
rect 34 -307007 50 -306973
rect -96 -307057 -62 -307041
rect -96 -308049 -62 -308033
rect 62 -307057 96 -307041
rect 62 -308049 96 -308033
rect -50 -308117 -34 -308083
rect 34 -308117 50 -308083
rect -50 -308225 -34 -308191
rect 34 -308225 50 -308191
rect -96 -308275 -62 -308259
rect -96 -309267 -62 -309251
rect 62 -308275 96 -308259
rect 62 -309267 96 -309251
rect -50 -309335 -34 -309301
rect 34 -309335 50 -309301
rect -50 -309443 -34 -309409
rect 34 -309443 50 -309409
rect -96 -309493 -62 -309477
rect -96 -310485 -62 -310469
rect 62 -309493 96 -309477
rect 62 -310485 96 -310469
rect -50 -310553 -34 -310519
rect 34 -310553 50 -310519
rect -50 -310661 -34 -310627
rect 34 -310661 50 -310627
rect -96 -310711 -62 -310695
rect -96 -311703 -62 -311687
rect 62 -310711 96 -310695
rect 62 -311703 96 -311687
rect -50 -311771 -34 -311737
rect 34 -311771 50 -311737
rect -50 -311879 -34 -311845
rect 34 -311879 50 -311845
rect -96 -311929 -62 -311913
rect -96 -312921 -62 -312905
rect 62 -311929 96 -311913
rect 62 -312921 96 -312905
rect -50 -312989 -34 -312955
rect 34 -312989 50 -312955
rect -50 -313097 -34 -313063
rect 34 -313097 50 -313063
rect -96 -313147 -62 -313131
rect -96 -314139 -62 -314123
rect 62 -313147 96 -313131
rect 62 -314139 96 -314123
rect -50 -314207 -34 -314173
rect 34 -314207 50 -314173
rect -50 -314315 -34 -314281
rect 34 -314315 50 -314281
rect -96 -314365 -62 -314349
rect -96 -315357 -62 -315341
rect 62 -314365 96 -314349
rect 62 -315357 96 -315341
rect -50 -315425 -34 -315391
rect 34 -315425 50 -315391
rect -50 -315533 -34 -315499
rect 34 -315533 50 -315499
rect -96 -315583 -62 -315567
rect -96 -316575 -62 -316559
rect 62 -315583 96 -315567
rect 62 -316575 96 -316559
rect -50 -316643 -34 -316609
rect 34 -316643 50 -316609
rect -50 -316751 -34 -316717
rect 34 -316751 50 -316717
rect -96 -316801 -62 -316785
rect -96 -317793 -62 -317777
rect 62 -316801 96 -316785
rect 62 -317793 96 -317777
rect -50 -317861 -34 -317827
rect 34 -317861 50 -317827
rect -50 -317969 -34 -317935
rect 34 -317969 50 -317935
rect -96 -318019 -62 -318003
rect -96 -319011 -62 -318995
rect 62 -318019 96 -318003
rect 62 -319011 96 -318995
rect -50 -319079 -34 -319045
rect 34 -319079 50 -319045
rect -50 -319187 -34 -319153
rect 34 -319187 50 -319153
rect -96 -319237 -62 -319221
rect -96 -320229 -62 -320213
rect 62 -319237 96 -319221
rect 62 -320229 96 -320213
rect -50 -320297 -34 -320263
rect 34 -320297 50 -320263
rect -50 -320405 -34 -320371
rect 34 -320405 50 -320371
rect -96 -320455 -62 -320439
rect -96 -321447 -62 -321431
rect 62 -320455 96 -320439
rect 62 -321447 96 -321431
rect -50 -321515 -34 -321481
rect 34 -321515 50 -321481
rect -50 -321623 -34 -321589
rect 34 -321623 50 -321589
rect -96 -321673 -62 -321657
rect -96 -322665 -62 -322649
rect 62 -321673 96 -321657
rect 62 -322665 96 -322649
rect -50 -322733 -34 -322699
rect 34 -322733 50 -322699
rect -50 -322841 -34 -322807
rect 34 -322841 50 -322807
rect -96 -322891 -62 -322875
rect -96 -323883 -62 -323867
rect 62 -322891 96 -322875
rect 62 -323883 96 -323867
rect -50 -323951 -34 -323917
rect 34 -323951 50 -323917
rect -50 -324059 -34 -324025
rect 34 -324059 50 -324025
rect -96 -324109 -62 -324093
rect -96 -325101 -62 -325085
rect 62 -324109 96 -324093
rect 62 -325101 96 -325085
rect -50 -325169 -34 -325135
rect 34 -325169 50 -325135
rect -50 -325277 -34 -325243
rect 34 -325277 50 -325243
rect -96 -325327 -62 -325311
rect -96 -326319 -62 -326303
rect 62 -325327 96 -325311
rect 62 -326319 96 -326303
rect -50 -326387 -34 -326353
rect 34 -326387 50 -326353
rect -50 -326495 -34 -326461
rect 34 -326495 50 -326461
rect -96 -326545 -62 -326529
rect -96 -327537 -62 -327521
rect 62 -326545 96 -326529
rect 62 -327537 96 -327521
rect -50 -327605 -34 -327571
rect 34 -327605 50 -327571
rect -50 -327713 -34 -327679
rect 34 -327713 50 -327679
rect -96 -327763 -62 -327747
rect -96 -328755 -62 -328739
rect 62 -327763 96 -327747
rect 62 -328755 96 -328739
rect -50 -328823 -34 -328789
rect 34 -328823 50 -328789
rect -50 -328931 -34 -328897
rect 34 -328931 50 -328897
rect -96 -328981 -62 -328965
rect -96 -329973 -62 -329957
rect 62 -328981 96 -328965
rect 62 -329973 96 -329957
rect -50 -330041 -34 -330007
rect 34 -330041 50 -330007
rect -50 -330149 -34 -330115
rect 34 -330149 50 -330115
rect -96 -330199 -62 -330183
rect -96 -331191 -62 -331175
rect 62 -330199 96 -330183
rect 62 -331191 96 -331175
rect -50 -331259 -34 -331225
rect 34 -331259 50 -331225
rect -50 -331367 -34 -331333
rect 34 -331367 50 -331333
rect -96 -331417 -62 -331401
rect -96 -332409 -62 -332393
rect 62 -331417 96 -331401
rect 62 -332409 96 -332393
rect -50 -332477 -34 -332443
rect 34 -332477 50 -332443
rect -50 -332585 -34 -332551
rect 34 -332585 50 -332551
rect -96 -332635 -62 -332619
rect -96 -333627 -62 -333611
rect 62 -332635 96 -332619
rect 62 -333627 96 -333611
rect -50 -333695 -34 -333661
rect 34 -333695 50 -333661
rect -50 -333803 -34 -333769
rect 34 -333803 50 -333769
rect -96 -333853 -62 -333837
rect -96 -334845 -62 -334829
rect 62 -333853 96 -333837
rect 62 -334845 96 -334829
rect -50 -334913 -34 -334879
rect 34 -334913 50 -334879
rect -50 -335021 -34 -334987
rect 34 -335021 50 -334987
rect -96 -335071 -62 -335055
rect -96 -336063 -62 -336047
rect 62 -335071 96 -335055
rect 62 -336063 96 -336047
rect -50 -336131 -34 -336097
rect 34 -336131 50 -336097
rect -50 -336239 -34 -336205
rect 34 -336239 50 -336205
rect -96 -336289 -62 -336273
rect -96 -337281 -62 -337265
rect 62 -336289 96 -336273
rect 62 -337281 96 -337265
rect -50 -337349 -34 -337315
rect 34 -337349 50 -337315
rect -50 -337457 -34 -337423
rect 34 -337457 50 -337423
rect -96 -337507 -62 -337491
rect -96 -338499 -62 -338483
rect 62 -337507 96 -337491
rect 62 -338499 96 -338483
rect -50 -338567 -34 -338533
rect 34 -338567 50 -338533
rect -50 -338675 -34 -338641
rect 34 -338675 50 -338641
rect -96 -338725 -62 -338709
rect -96 -339717 -62 -339701
rect 62 -338725 96 -338709
rect 62 -339717 96 -339701
rect -50 -339785 -34 -339751
rect 34 -339785 50 -339751
rect -50 -339893 -34 -339859
rect 34 -339893 50 -339859
rect -96 -339943 -62 -339927
rect -96 -340935 -62 -340919
rect 62 -339943 96 -339927
rect 62 -340935 96 -340919
rect -50 -341003 -34 -340969
rect 34 -341003 50 -340969
rect -50 -341111 -34 -341077
rect 34 -341111 50 -341077
rect -96 -341161 -62 -341145
rect -96 -342153 -62 -342137
rect 62 -341161 96 -341145
rect 62 -342153 96 -342137
rect -50 -342221 -34 -342187
rect 34 -342221 50 -342187
rect -50 -342329 -34 -342295
rect 34 -342329 50 -342295
rect -96 -342379 -62 -342363
rect -96 -343371 -62 -343355
rect 62 -342379 96 -342363
rect 62 -343371 96 -343355
rect -50 -343439 -34 -343405
rect 34 -343439 50 -343405
rect -50 -343547 -34 -343513
rect 34 -343547 50 -343513
rect -96 -343597 -62 -343581
rect -96 -344589 -62 -344573
rect 62 -343597 96 -343581
rect 62 -344589 96 -344573
rect -50 -344657 -34 -344623
rect 34 -344657 50 -344623
rect -50 -344765 -34 -344731
rect 34 -344765 50 -344731
rect -96 -344815 -62 -344799
rect -96 -345807 -62 -345791
rect 62 -344815 96 -344799
rect 62 -345807 96 -345791
rect -50 -345875 -34 -345841
rect 34 -345875 50 -345841
rect -50 -345983 -34 -345949
rect 34 -345983 50 -345949
rect -96 -346033 -62 -346017
rect -96 -347025 -62 -347009
rect 62 -346033 96 -346017
rect 62 -347025 96 -347009
rect -50 -347093 -34 -347059
rect 34 -347093 50 -347059
rect -50 -347201 -34 -347167
rect 34 -347201 50 -347167
rect -96 -347251 -62 -347235
rect -96 -348243 -62 -348227
rect 62 -347251 96 -347235
rect 62 -348243 96 -348227
rect -50 -348311 -34 -348277
rect 34 -348311 50 -348277
rect -50 -348419 -34 -348385
rect 34 -348419 50 -348385
rect -96 -348469 -62 -348453
rect -96 -349461 -62 -349445
rect 62 -348469 96 -348453
rect 62 -349461 96 -349445
rect -50 -349529 -34 -349495
rect 34 -349529 50 -349495
rect -50 -349637 -34 -349603
rect 34 -349637 50 -349603
rect -96 -349687 -62 -349671
rect -96 -350679 -62 -350663
rect 62 -349687 96 -349671
rect 62 -350679 96 -350663
rect -50 -350747 -34 -350713
rect 34 -350747 50 -350713
rect -50 -350855 -34 -350821
rect 34 -350855 50 -350821
rect -96 -350905 -62 -350889
rect -96 -351897 -62 -351881
rect 62 -350905 96 -350889
rect 62 -351897 96 -351881
rect -50 -351965 -34 -351931
rect 34 -351965 50 -351931
rect -50 -352073 -34 -352039
rect 34 -352073 50 -352039
rect -96 -352123 -62 -352107
rect -96 -353115 -62 -353099
rect 62 -352123 96 -352107
rect 62 -353115 96 -353099
rect -50 -353183 -34 -353149
rect 34 -353183 50 -353149
rect -50 -353291 -34 -353257
rect 34 -353291 50 -353257
rect -96 -353341 -62 -353325
rect -96 -354333 -62 -354317
rect 62 -353341 96 -353325
rect 62 -354333 96 -354317
rect -50 -354401 -34 -354367
rect 34 -354401 50 -354367
rect -50 -354509 -34 -354475
rect 34 -354509 50 -354475
rect -96 -354559 -62 -354543
rect -96 -355551 -62 -355535
rect 62 -354559 96 -354543
rect 62 -355551 96 -355535
rect -50 -355619 -34 -355585
rect 34 -355619 50 -355585
rect -50 -355727 -34 -355693
rect 34 -355727 50 -355693
rect -96 -355777 -62 -355761
rect -96 -356769 -62 -356753
rect 62 -355777 96 -355761
rect 62 -356769 96 -356753
rect -50 -356837 -34 -356803
rect 34 -356837 50 -356803
rect -50 -356945 -34 -356911
rect 34 -356945 50 -356911
rect -96 -356995 -62 -356979
rect -96 -357987 -62 -357971
rect 62 -356995 96 -356979
rect 62 -357987 96 -357971
rect -50 -358055 -34 -358021
rect 34 -358055 50 -358021
rect -50 -358163 -34 -358129
rect 34 -358163 50 -358129
rect -96 -358213 -62 -358197
rect -96 -359205 -62 -359189
rect 62 -358213 96 -358197
rect 62 -359205 96 -359189
rect -50 -359273 -34 -359239
rect 34 -359273 50 -359239
rect -50 -359381 -34 -359347
rect 34 -359381 50 -359347
rect -96 -359431 -62 -359415
rect -96 -360423 -62 -360407
rect 62 -359431 96 -359415
rect 62 -360423 96 -360407
rect -50 -360491 -34 -360457
rect 34 -360491 50 -360457
rect -50 -360599 -34 -360565
rect 34 -360599 50 -360565
rect -96 -360649 -62 -360633
rect -96 -361641 -62 -361625
rect 62 -360649 96 -360633
rect 62 -361641 96 -361625
rect -50 -361709 -34 -361675
rect 34 -361709 50 -361675
rect -50 -361817 -34 -361783
rect 34 -361817 50 -361783
rect -96 -361867 -62 -361851
rect -96 -362859 -62 -362843
rect 62 -361867 96 -361851
rect 62 -362859 96 -362843
rect -50 -362927 -34 -362893
rect 34 -362927 50 -362893
rect -50 -363035 -34 -363001
rect 34 -363035 50 -363001
rect -96 -363085 -62 -363069
rect -96 -364077 -62 -364061
rect 62 -363085 96 -363069
rect 62 -364077 96 -364061
rect -50 -364145 -34 -364111
rect 34 -364145 50 -364111
rect -50 -364253 -34 -364219
rect 34 -364253 50 -364219
rect -96 -364303 -62 -364287
rect -96 -365295 -62 -365279
rect 62 -364303 96 -364287
rect 62 -365295 96 -365279
rect -50 -365363 -34 -365329
rect 34 -365363 50 -365329
rect -50 -365471 -34 -365437
rect 34 -365471 50 -365437
rect -96 -365521 -62 -365505
rect -96 -366513 -62 -366497
rect 62 -365521 96 -365505
rect 62 -366513 96 -366497
rect -50 -366581 -34 -366547
rect 34 -366581 50 -366547
rect -50 -366689 -34 -366655
rect 34 -366689 50 -366655
rect -96 -366739 -62 -366723
rect -96 -367731 -62 -367715
rect 62 -366739 96 -366723
rect 62 -367731 96 -367715
rect -50 -367799 -34 -367765
rect 34 -367799 50 -367765
rect -50 -367907 -34 -367873
rect 34 -367907 50 -367873
rect -96 -367957 -62 -367941
rect -96 -368949 -62 -368933
rect 62 -367957 96 -367941
rect 62 -368949 96 -368933
rect -50 -369017 -34 -368983
rect 34 -369017 50 -368983
rect -50 -369125 -34 -369091
rect 34 -369125 50 -369091
rect -96 -369175 -62 -369159
rect -96 -370167 -62 -370151
rect 62 -369175 96 -369159
rect 62 -370167 96 -370151
rect -50 -370235 -34 -370201
rect 34 -370235 50 -370201
rect -50 -370343 -34 -370309
rect 34 -370343 50 -370309
rect -96 -370393 -62 -370377
rect -96 -371385 -62 -371369
rect 62 -370393 96 -370377
rect 62 -371385 96 -371369
rect -50 -371453 -34 -371419
rect 34 -371453 50 -371419
rect -50 -371561 -34 -371527
rect 34 -371561 50 -371527
rect -96 -371611 -62 -371595
rect -96 -372603 -62 -372587
rect 62 -371611 96 -371595
rect 62 -372603 96 -372587
rect -50 -372671 -34 -372637
rect 34 -372671 50 -372637
rect -50 -372779 -34 -372745
rect 34 -372779 50 -372745
rect -96 -372829 -62 -372813
rect -96 -373821 -62 -373805
rect 62 -372829 96 -372813
rect 62 -373821 96 -373805
rect -50 -373889 -34 -373855
rect 34 -373889 50 -373855
rect -50 -373997 -34 -373963
rect 34 -373997 50 -373963
rect -96 -374047 -62 -374031
rect -96 -375039 -62 -375023
rect 62 -374047 96 -374031
rect 62 -375039 96 -375023
rect -50 -375107 -34 -375073
rect 34 -375107 50 -375073
rect -50 -375215 -34 -375181
rect 34 -375215 50 -375181
rect -96 -375265 -62 -375249
rect -96 -376257 -62 -376241
rect 62 -375265 96 -375249
rect 62 -376257 96 -376241
rect -50 -376325 -34 -376291
rect 34 -376325 50 -376291
rect -50 -376433 -34 -376399
rect 34 -376433 50 -376399
rect -96 -376483 -62 -376467
rect -96 -377475 -62 -377459
rect 62 -376483 96 -376467
rect 62 -377475 96 -377459
rect -50 -377543 -34 -377509
rect 34 -377543 50 -377509
rect -50 -377651 -34 -377617
rect 34 -377651 50 -377617
rect -96 -377701 -62 -377685
rect -96 -378693 -62 -378677
rect 62 -377701 96 -377685
rect 62 -378693 96 -378677
rect -50 -378761 -34 -378727
rect 34 -378761 50 -378727
rect -50 -378869 -34 -378835
rect 34 -378869 50 -378835
rect -96 -378919 -62 -378903
rect -96 -379911 -62 -379895
rect 62 -378919 96 -378903
rect 62 -379911 96 -379895
rect -50 -379979 -34 -379945
rect 34 -379979 50 -379945
rect -50 -380087 -34 -380053
rect 34 -380087 50 -380053
rect -96 -380137 -62 -380121
rect -96 -381129 -62 -381113
rect 62 -380137 96 -380121
rect 62 -381129 96 -381113
rect -50 -381197 -34 -381163
rect 34 -381197 50 -381163
rect -50 -381305 -34 -381271
rect 34 -381305 50 -381271
rect -96 -381355 -62 -381339
rect -96 -382347 -62 -382331
rect 62 -381355 96 -381339
rect 62 -382347 96 -382331
rect -50 -382415 -34 -382381
rect 34 -382415 50 -382381
rect -50 -382523 -34 -382489
rect 34 -382523 50 -382489
rect -96 -382573 -62 -382557
rect -96 -383565 -62 -383549
rect 62 -382573 96 -382557
rect 62 -383565 96 -383549
rect -50 -383633 -34 -383599
rect 34 -383633 50 -383599
rect -50 -383741 -34 -383707
rect 34 -383741 50 -383707
rect -96 -383791 -62 -383775
rect -96 -384783 -62 -384767
rect 62 -383791 96 -383775
rect 62 -384783 96 -384767
rect -50 -384851 -34 -384817
rect 34 -384851 50 -384817
rect -50 -384959 -34 -384925
rect 34 -384959 50 -384925
rect -96 -385009 -62 -384993
rect -96 -386001 -62 -385985
rect 62 -385009 96 -384993
rect 62 -386001 96 -385985
rect -50 -386069 -34 -386035
rect 34 -386069 50 -386035
rect -50 -386177 -34 -386143
rect 34 -386177 50 -386143
rect -96 -386227 -62 -386211
rect -96 -387219 -62 -387203
rect 62 -386227 96 -386211
rect 62 -387219 96 -387203
rect -50 -387287 -34 -387253
rect 34 -387287 50 -387253
rect -50 -387395 -34 -387361
rect 34 -387395 50 -387361
rect -96 -387445 -62 -387429
rect -96 -388437 -62 -388421
rect 62 -387445 96 -387429
rect 62 -388437 96 -388421
rect -50 -388505 -34 -388471
rect 34 -388505 50 -388471
rect -50 -388613 -34 -388579
rect 34 -388613 50 -388579
rect -96 -388663 -62 -388647
rect -96 -389655 -62 -389639
rect 62 -388663 96 -388647
rect 62 -389655 96 -389639
rect -50 -389723 -34 -389689
rect 34 -389723 50 -389689
rect -50 -389831 -34 -389797
rect 34 -389831 50 -389797
rect -96 -389881 -62 -389865
rect -96 -390873 -62 -390857
rect 62 -389881 96 -389865
rect 62 -390873 96 -390857
rect -50 -390941 -34 -390907
rect 34 -390941 50 -390907
rect -50 -391049 -34 -391015
rect 34 -391049 50 -391015
rect -96 -391099 -62 -391083
rect -96 -392091 -62 -392075
rect 62 -391099 96 -391083
rect 62 -392091 96 -392075
rect -50 -392159 -34 -392125
rect 34 -392159 50 -392125
rect -50 -392267 -34 -392233
rect 34 -392267 50 -392233
rect -96 -392317 -62 -392301
rect -96 -393309 -62 -393293
rect 62 -392317 96 -392301
rect 62 -393309 96 -393293
rect -50 -393377 -34 -393343
rect 34 -393377 50 -393343
rect -50 -393485 -34 -393451
rect 34 -393485 50 -393451
rect -96 -393535 -62 -393519
rect -96 -394527 -62 -394511
rect 62 -393535 96 -393519
rect 62 -394527 96 -394511
rect -50 -394595 -34 -394561
rect 34 -394595 50 -394561
rect -50 -394703 -34 -394669
rect 34 -394703 50 -394669
rect -96 -394753 -62 -394737
rect -96 -395745 -62 -395729
rect 62 -394753 96 -394737
rect 62 -395745 96 -395729
rect -50 -395813 -34 -395779
rect 34 -395813 50 -395779
rect -50 -395921 -34 -395887
rect 34 -395921 50 -395887
rect -96 -395971 -62 -395955
rect -96 -396963 -62 -396947
rect 62 -395971 96 -395955
rect 62 -396963 96 -396947
rect -50 -397031 -34 -396997
rect 34 -397031 50 -396997
rect -50 -397139 -34 -397105
rect 34 -397139 50 -397105
rect -96 -397189 -62 -397173
rect -96 -398181 -62 -398165
rect 62 -397189 96 -397173
rect 62 -398181 96 -398165
rect -50 -398249 -34 -398215
rect 34 -398249 50 -398215
rect -50 -398357 -34 -398323
rect 34 -398357 50 -398323
rect -96 -398407 -62 -398391
rect -96 -399399 -62 -399383
rect 62 -398407 96 -398391
rect 62 -399399 96 -399383
rect -50 -399467 -34 -399433
rect 34 -399467 50 -399433
rect -50 -399575 -34 -399541
rect 34 -399575 50 -399541
rect -96 -399625 -62 -399609
rect -96 -400617 -62 -400601
rect 62 -399625 96 -399609
rect 62 -400617 96 -400601
rect -50 -400685 -34 -400651
rect 34 -400685 50 -400651
rect -50 -400793 -34 -400759
rect 34 -400793 50 -400759
rect -96 -400843 -62 -400827
rect -96 -401835 -62 -401819
rect 62 -400843 96 -400827
rect 62 -401835 96 -401819
rect -50 -401903 -34 -401869
rect 34 -401903 50 -401869
rect -50 -402011 -34 -401977
rect 34 -402011 50 -401977
rect -96 -402061 -62 -402045
rect -96 -403053 -62 -403037
rect 62 -402061 96 -402045
rect 62 -403053 96 -403037
rect -50 -403121 -34 -403087
rect 34 -403121 50 -403087
rect -50 -403229 -34 -403195
rect 34 -403229 50 -403195
rect -96 -403279 -62 -403263
rect -96 -404271 -62 -404255
rect 62 -403279 96 -403263
rect 62 -404271 96 -404255
rect -50 -404339 -34 -404305
rect 34 -404339 50 -404305
rect -50 -404447 -34 -404413
rect 34 -404447 50 -404413
rect -96 -404497 -62 -404481
rect -96 -405489 -62 -405473
rect 62 -404497 96 -404481
rect 62 -405489 96 -405473
rect -50 -405557 -34 -405523
rect 34 -405557 50 -405523
rect -50 -405665 -34 -405631
rect 34 -405665 50 -405631
rect -96 -405715 -62 -405699
rect -96 -406707 -62 -406691
rect 62 -405715 96 -405699
rect 62 -406707 96 -406691
rect -50 -406775 -34 -406741
rect 34 -406775 50 -406741
rect -50 -406883 -34 -406849
rect 34 -406883 50 -406849
rect -96 -406933 -62 -406917
rect -96 -407925 -62 -407909
rect 62 -406933 96 -406917
rect 62 -407925 96 -407909
rect -50 -407993 -34 -407959
rect 34 -407993 50 -407959
rect -50 -408101 -34 -408067
rect 34 -408101 50 -408067
rect -96 -408151 -62 -408135
rect -96 -409143 -62 -409127
rect 62 -408151 96 -408135
rect 62 -409143 96 -409127
rect -50 -409211 -34 -409177
rect 34 -409211 50 -409177
rect -50 -409319 -34 -409285
rect 34 -409319 50 -409285
rect -96 -409369 -62 -409353
rect -96 -410361 -62 -410345
rect 62 -409369 96 -409353
rect 62 -410361 96 -410345
rect -50 -410429 -34 -410395
rect 34 -410429 50 -410395
rect -50 -410537 -34 -410503
rect 34 -410537 50 -410503
rect -96 -410587 -62 -410571
rect -96 -411579 -62 -411563
rect 62 -410587 96 -410571
rect 62 -411579 96 -411563
rect -50 -411647 -34 -411613
rect 34 -411647 50 -411613
rect -50 -411755 -34 -411721
rect 34 -411755 50 -411721
rect -96 -411805 -62 -411789
rect -96 -412797 -62 -412781
rect 62 -411805 96 -411789
rect 62 -412797 96 -412781
rect -50 -412865 -34 -412831
rect 34 -412865 50 -412831
rect -50 -412973 -34 -412939
rect 34 -412973 50 -412939
rect -96 -413023 -62 -413007
rect -96 -414015 -62 -413999
rect 62 -413023 96 -413007
rect 62 -414015 96 -413999
rect -50 -414083 -34 -414049
rect 34 -414083 50 -414049
rect -50 -414191 -34 -414157
rect 34 -414191 50 -414157
rect -96 -414241 -62 -414225
rect -96 -415233 -62 -415217
rect 62 -414241 96 -414225
rect 62 -415233 96 -415217
rect -50 -415301 -34 -415267
rect 34 -415301 50 -415267
rect -50 -415409 -34 -415375
rect 34 -415409 50 -415375
rect -96 -415459 -62 -415443
rect -96 -416451 -62 -416435
rect 62 -415459 96 -415443
rect 62 -416451 96 -416435
rect -50 -416519 -34 -416485
rect 34 -416519 50 -416485
rect -50 -416627 -34 -416593
rect 34 -416627 50 -416593
rect -96 -416677 -62 -416661
rect -96 -417669 -62 -417653
rect 62 -416677 96 -416661
rect 62 -417669 96 -417653
rect -50 -417737 -34 -417703
rect 34 -417737 50 -417703
rect -50 -417845 -34 -417811
rect 34 -417845 50 -417811
rect -96 -417895 -62 -417879
rect -96 -418887 -62 -418871
rect 62 -417895 96 -417879
rect 62 -418887 96 -418871
rect -50 -418955 -34 -418921
rect 34 -418955 50 -418921
rect -50 -419063 -34 -419029
rect 34 -419063 50 -419029
rect -96 -419113 -62 -419097
rect -96 -420105 -62 -420089
rect 62 -419113 96 -419097
rect 62 -420105 96 -420089
rect -50 -420173 -34 -420139
rect 34 -420173 50 -420139
rect -50 -420281 -34 -420247
rect 34 -420281 50 -420247
rect -96 -420331 -62 -420315
rect -96 -421323 -62 -421307
rect 62 -420331 96 -420315
rect 62 -421323 96 -421307
rect -50 -421391 -34 -421357
rect 34 -421391 50 -421357
rect -50 -421499 -34 -421465
rect 34 -421499 50 -421465
rect -96 -421549 -62 -421533
rect -96 -422541 -62 -422525
rect 62 -421549 96 -421533
rect 62 -422541 96 -422525
rect -50 -422609 -34 -422575
rect 34 -422609 50 -422575
rect -50 -422717 -34 -422683
rect 34 -422717 50 -422683
rect -96 -422767 -62 -422751
rect -96 -423759 -62 -423743
rect 62 -422767 96 -422751
rect 62 -423759 96 -423743
rect -50 -423827 -34 -423793
rect 34 -423827 50 -423793
rect -50 -423935 -34 -423901
rect 34 -423935 50 -423901
rect -96 -423985 -62 -423969
rect -96 -424977 -62 -424961
rect 62 -423985 96 -423969
rect 62 -424977 96 -424961
rect -50 -425045 -34 -425011
rect 34 -425045 50 -425011
rect -50 -425153 -34 -425119
rect 34 -425153 50 -425119
rect -96 -425203 -62 -425187
rect -96 -426195 -62 -426179
rect 62 -425203 96 -425187
rect 62 -426195 96 -426179
rect -50 -426263 -34 -426229
rect 34 -426263 50 -426229
rect -50 -426371 -34 -426337
rect 34 -426371 50 -426337
rect -96 -426421 -62 -426405
rect -96 -427413 -62 -427397
rect 62 -426421 96 -426405
rect 62 -427413 96 -427397
rect -50 -427481 -34 -427447
rect 34 -427481 50 -427447
rect -50 -427589 -34 -427555
rect 34 -427589 50 -427555
rect -96 -427639 -62 -427623
rect -96 -428631 -62 -428615
rect 62 -427639 96 -427623
rect 62 -428631 96 -428615
rect -50 -428699 -34 -428665
rect 34 -428699 50 -428665
rect -50 -428807 -34 -428773
rect 34 -428807 50 -428773
rect -96 -428857 -62 -428841
rect -96 -429849 -62 -429833
rect 62 -428857 96 -428841
rect 62 -429849 96 -429833
rect -50 -429917 -34 -429883
rect 34 -429917 50 -429883
rect -50 -430025 -34 -429991
rect 34 -430025 50 -429991
rect -96 -430075 -62 -430059
rect -96 -431067 -62 -431051
rect 62 -430075 96 -430059
rect 62 -431067 96 -431051
rect -50 -431135 -34 -431101
rect 34 -431135 50 -431101
rect -50 -431243 -34 -431209
rect 34 -431243 50 -431209
rect -96 -431293 -62 -431277
rect -96 -432285 -62 -432269
rect 62 -431293 96 -431277
rect 62 -432285 96 -432269
rect -50 -432353 -34 -432319
rect 34 -432353 50 -432319
rect -50 -432461 -34 -432427
rect 34 -432461 50 -432427
rect -96 -432511 -62 -432495
rect -96 -433503 -62 -433487
rect 62 -432511 96 -432495
rect 62 -433503 96 -433487
rect -50 -433571 -34 -433537
rect 34 -433571 50 -433537
rect -50 -433679 -34 -433645
rect 34 -433679 50 -433645
rect -96 -433729 -62 -433713
rect -96 -434721 -62 -434705
rect 62 -433729 96 -433713
rect 62 -434721 96 -434705
rect -50 -434789 -34 -434755
rect 34 -434789 50 -434755
rect -50 -434897 -34 -434863
rect 34 -434897 50 -434863
rect -96 -434947 -62 -434931
rect -96 -435939 -62 -435923
rect 62 -434947 96 -434931
rect 62 -435939 96 -435923
rect -50 -436007 -34 -435973
rect 34 -436007 50 -435973
rect -50 -436115 -34 -436081
rect 34 -436115 50 -436081
rect -96 -436165 -62 -436149
rect -96 -437157 -62 -437141
rect 62 -436165 96 -436149
rect 62 -437157 96 -437141
rect -50 -437225 -34 -437191
rect 34 -437225 50 -437191
rect -50 -437333 -34 -437299
rect 34 -437333 50 -437299
rect -96 -437383 -62 -437367
rect -96 -438375 -62 -438359
rect 62 -437383 96 -437367
rect 62 -438375 96 -438359
rect -50 -438443 -34 -438409
rect 34 -438443 50 -438409
rect -50 -438551 -34 -438517
rect 34 -438551 50 -438517
rect -96 -438601 -62 -438585
rect -96 -439593 -62 -439577
rect 62 -438601 96 -438585
rect 62 -439593 96 -439577
rect -50 -439661 -34 -439627
rect 34 -439661 50 -439627
rect -50 -439769 -34 -439735
rect 34 -439769 50 -439735
rect -96 -439819 -62 -439803
rect -96 -440811 -62 -440795
rect 62 -439819 96 -439803
rect 62 -440811 96 -440795
rect -50 -440879 -34 -440845
rect 34 -440879 50 -440845
rect -50 -440987 -34 -440953
rect 34 -440987 50 -440953
rect -96 -441037 -62 -441021
rect -96 -442029 -62 -442013
rect 62 -441037 96 -441021
rect 62 -442029 96 -442013
rect -50 -442097 -34 -442063
rect 34 -442097 50 -442063
rect -50 -442205 -34 -442171
rect 34 -442205 50 -442171
rect -96 -442255 -62 -442239
rect -96 -443247 -62 -443231
rect 62 -442255 96 -442239
rect 62 -443247 96 -443231
rect -50 -443315 -34 -443281
rect 34 -443315 50 -443281
rect -50 -443423 -34 -443389
rect 34 -443423 50 -443389
rect -96 -443473 -62 -443457
rect -96 -444465 -62 -444449
rect 62 -443473 96 -443457
rect 62 -444465 96 -444449
rect -50 -444533 -34 -444499
rect 34 -444533 50 -444499
rect -50 -444641 -34 -444607
rect 34 -444641 50 -444607
rect -96 -444691 -62 -444675
rect -96 -445683 -62 -445667
rect 62 -444691 96 -444675
rect 62 -445683 96 -445667
rect -50 -445751 -34 -445717
rect 34 -445751 50 -445717
rect -50 -445859 -34 -445825
rect 34 -445859 50 -445825
rect -96 -445909 -62 -445893
rect -96 -446901 -62 -446885
rect 62 -445909 96 -445893
rect 62 -446901 96 -446885
rect -50 -446969 -34 -446935
rect 34 -446969 50 -446935
rect -50 -447077 -34 -447043
rect 34 -447077 50 -447043
rect -96 -447127 -62 -447111
rect -96 -448119 -62 -448103
rect 62 -447127 96 -447111
rect 62 -448119 96 -448103
rect -50 -448187 -34 -448153
rect 34 -448187 50 -448153
rect -50 -448295 -34 -448261
rect 34 -448295 50 -448261
rect -96 -448345 -62 -448329
rect -96 -449337 -62 -449321
rect 62 -448345 96 -448329
rect 62 -449337 96 -449321
rect -50 -449405 -34 -449371
rect 34 -449405 50 -449371
rect -50 -449513 -34 -449479
rect 34 -449513 50 -449479
rect -96 -449563 -62 -449547
rect -96 -450555 -62 -450539
rect 62 -449563 96 -449547
rect 62 -450555 96 -450539
rect -50 -450623 -34 -450589
rect 34 -450623 50 -450589
rect -50 -450731 -34 -450697
rect 34 -450731 50 -450697
rect -96 -450781 -62 -450765
rect -96 -451773 -62 -451757
rect 62 -450781 96 -450765
rect 62 -451773 96 -451757
rect -50 -451841 -34 -451807
rect 34 -451841 50 -451807
rect -50 -451949 -34 -451915
rect 34 -451949 50 -451915
rect -96 -451999 -62 -451983
rect -96 -452991 -62 -452975
rect 62 -451999 96 -451983
rect 62 -452991 96 -452975
rect -50 -453059 -34 -453025
rect 34 -453059 50 -453025
rect -50 -453167 -34 -453133
rect 34 -453167 50 -453133
rect -96 -453217 -62 -453201
rect -96 -454209 -62 -454193
rect 62 -453217 96 -453201
rect 62 -454209 96 -454193
rect -50 -454277 -34 -454243
rect 34 -454277 50 -454243
rect -50 -454385 -34 -454351
rect 34 -454385 50 -454351
rect -96 -454435 -62 -454419
rect -96 -455427 -62 -455411
rect 62 -454435 96 -454419
rect 62 -455427 96 -455411
rect -50 -455495 -34 -455461
rect 34 -455495 50 -455461
rect -50 -455603 -34 -455569
rect 34 -455603 50 -455569
rect -96 -455653 -62 -455637
rect -96 -456645 -62 -456629
rect 62 -455653 96 -455637
rect 62 -456645 96 -456629
rect -50 -456713 -34 -456679
rect 34 -456713 50 -456679
rect -50 -456821 -34 -456787
rect 34 -456821 50 -456787
rect -96 -456871 -62 -456855
rect -96 -457863 -62 -457847
rect 62 -456871 96 -456855
rect 62 -457863 96 -457847
rect -50 -457931 -34 -457897
rect 34 -457931 50 -457897
rect -50 -458039 -34 -458005
rect 34 -458039 50 -458005
rect -96 -458089 -62 -458073
rect -96 -459081 -62 -459065
rect 62 -458089 96 -458073
rect 62 -459081 96 -459065
rect -50 -459149 -34 -459115
rect 34 -459149 50 -459115
rect -50 -459257 -34 -459223
rect 34 -459257 50 -459223
rect -96 -459307 -62 -459291
rect -96 -460299 -62 -460283
rect 62 -459307 96 -459291
rect 62 -460299 96 -460283
rect -50 -460367 -34 -460333
rect 34 -460367 50 -460333
rect -50 -460475 -34 -460441
rect 34 -460475 50 -460441
rect -96 -460525 -62 -460509
rect -96 -461517 -62 -461501
rect 62 -460525 96 -460509
rect 62 -461517 96 -461501
rect -50 -461585 -34 -461551
rect 34 -461585 50 -461551
rect -50 -461693 -34 -461659
rect 34 -461693 50 -461659
rect -96 -461743 -62 -461727
rect -96 -462735 -62 -462719
rect 62 -461743 96 -461727
rect 62 -462735 96 -462719
rect -50 -462803 -34 -462769
rect 34 -462803 50 -462769
rect -50 -462911 -34 -462877
rect 34 -462911 50 -462877
rect -96 -462961 -62 -462945
rect -96 -463953 -62 -463937
rect 62 -462961 96 -462945
rect 62 -463953 96 -463937
rect -50 -464021 -34 -463987
rect 34 -464021 50 -463987
rect -50 -464129 -34 -464095
rect 34 -464129 50 -464095
rect -96 -464179 -62 -464163
rect -96 -465171 -62 -465155
rect 62 -464179 96 -464163
rect 62 -465171 96 -465155
rect -50 -465239 -34 -465205
rect 34 -465239 50 -465205
rect -50 -465347 -34 -465313
rect 34 -465347 50 -465313
rect -96 -465397 -62 -465381
rect -96 -466389 -62 -466373
rect 62 -465397 96 -465381
rect 62 -466389 96 -466373
rect -50 -466457 -34 -466423
rect 34 -466457 50 -466423
rect -50 -466565 -34 -466531
rect 34 -466565 50 -466531
rect -96 -466615 -62 -466599
rect -96 -467607 -62 -467591
rect 62 -466615 96 -466599
rect 62 -467607 96 -467591
rect -50 -467675 -34 -467641
rect 34 -467675 50 -467641
rect -50 -467783 -34 -467749
rect 34 -467783 50 -467749
rect -96 -467833 -62 -467817
rect -96 -468825 -62 -468809
rect 62 -467833 96 -467817
rect 62 -468825 96 -468809
rect -50 -468893 -34 -468859
rect 34 -468893 50 -468859
rect -50 -469001 -34 -468967
rect 34 -469001 50 -468967
rect -96 -469051 -62 -469035
rect -96 -470043 -62 -470027
rect 62 -469051 96 -469035
rect 62 -470043 96 -470027
rect -50 -470111 -34 -470077
rect 34 -470111 50 -470077
rect -50 -470219 -34 -470185
rect 34 -470219 50 -470185
rect -96 -470269 -62 -470253
rect -96 -471261 -62 -471245
rect 62 -470269 96 -470253
rect 62 -471261 96 -471245
rect -50 -471329 -34 -471295
rect 34 -471329 50 -471295
rect -50 -471437 -34 -471403
rect 34 -471437 50 -471403
rect -96 -471487 -62 -471471
rect -96 -472479 -62 -472463
rect 62 -471487 96 -471471
rect 62 -472479 96 -472463
rect -50 -472547 -34 -472513
rect 34 -472547 50 -472513
rect -50 -472655 -34 -472621
rect 34 -472655 50 -472621
rect -96 -472705 -62 -472689
rect -96 -473697 -62 -473681
rect 62 -472705 96 -472689
rect 62 -473697 96 -473681
rect -50 -473765 -34 -473731
rect 34 -473765 50 -473731
rect -50 -473873 -34 -473839
rect 34 -473873 50 -473839
rect -96 -473923 -62 -473907
rect -96 -474915 -62 -474899
rect 62 -473923 96 -473907
rect 62 -474915 96 -474899
rect -50 -474983 -34 -474949
rect 34 -474983 50 -474949
rect -50 -475091 -34 -475057
rect 34 -475091 50 -475057
rect -96 -475141 -62 -475125
rect -96 -476133 -62 -476117
rect 62 -475141 96 -475125
rect 62 -476133 96 -476117
rect -50 -476201 -34 -476167
rect 34 -476201 50 -476167
rect -50 -476309 -34 -476275
rect 34 -476309 50 -476275
rect -96 -476359 -62 -476343
rect -96 -477351 -62 -477335
rect 62 -476359 96 -476343
rect 62 -477351 96 -477335
rect -50 -477419 -34 -477385
rect 34 -477419 50 -477385
rect -50 -477527 -34 -477493
rect 34 -477527 50 -477493
rect -96 -477577 -62 -477561
rect -96 -478569 -62 -478553
rect 62 -477577 96 -477561
rect 62 -478569 96 -478553
rect -50 -478637 -34 -478603
rect 34 -478637 50 -478603
rect -50 -478745 -34 -478711
rect 34 -478745 50 -478711
rect -96 -478795 -62 -478779
rect -96 -479787 -62 -479771
rect 62 -478795 96 -478779
rect 62 -479787 96 -479771
rect -50 -479855 -34 -479821
rect 34 -479855 50 -479821
rect -50 -479963 -34 -479929
rect 34 -479963 50 -479929
rect -96 -480013 -62 -479997
rect -96 -481005 -62 -480989
rect 62 -480013 96 -479997
rect 62 -481005 96 -480989
rect -50 -481073 -34 -481039
rect 34 -481073 50 -481039
rect -50 -481181 -34 -481147
rect 34 -481181 50 -481147
rect -96 -481231 -62 -481215
rect -96 -482223 -62 -482207
rect 62 -481231 96 -481215
rect 62 -482223 96 -482207
rect -50 -482291 -34 -482257
rect 34 -482291 50 -482257
rect -50 -482399 -34 -482365
rect 34 -482399 50 -482365
rect -96 -482449 -62 -482433
rect -96 -483441 -62 -483425
rect 62 -482449 96 -482433
rect 62 -483441 96 -483425
rect -50 -483509 -34 -483475
rect 34 -483509 50 -483475
rect -50 -483617 -34 -483583
rect 34 -483617 50 -483583
rect -96 -483667 -62 -483651
rect -96 -484659 -62 -484643
rect 62 -483667 96 -483651
rect 62 -484659 96 -484643
rect -50 -484727 -34 -484693
rect 34 -484727 50 -484693
rect -50 -484835 -34 -484801
rect 34 -484835 50 -484801
rect -96 -484885 -62 -484869
rect -96 -485877 -62 -485861
rect 62 -484885 96 -484869
rect 62 -485877 96 -485861
rect -50 -485945 -34 -485911
rect 34 -485945 50 -485911
rect -50 -486053 -34 -486019
rect 34 -486053 50 -486019
rect -96 -486103 -62 -486087
rect -96 -487095 -62 -487079
rect 62 -486103 96 -486087
rect 62 -487095 96 -487079
rect -50 -487163 -34 -487129
rect 34 -487163 50 -487129
rect -50 -487271 -34 -487237
rect 34 -487271 50 -487237
rect -96 -487321 -62 -487305
rect -96 -488313 -62 -488297
rect 62 -487321 96 -487305
rect 62 -488313 96 -488297
rect -50 -488381 -34 -488347
rect 34 -488381 50 -488347
rect -50 -488489 -34 -488455
rect 34 -488489 50 -488455
rect -96 -488539 -62 -488523
rect -96 -489531 -62 -489515
rect 62 -488539 96 -488523
rect 62 -489531 96 -489515
rect -50 -489599 -34 -489565
rect 34 -489599 50 -489565
rect -50 -489707 -34 -489673
rect 34 -489707 50 -489673
rect -96 -489757 -62 -489741
rect -96 -490749 -62 -490733
rect 62 -489757 96 -489741
rect 62 -490749 96 -490733
rect -50 -490817 -34 -490783
rect 34 -490817 50 -490783
rect -50 -490925 -34 -490891
rect 34 -490925 50 -490891
rect -96 -490975 -62 -490959
rect -96 -491967 -62 -491951
rect 62 -490975 96 -490959
rect 62 -491967 96 -491951
rect -50 -492035 -34 -492001
rect 34 -492035 50 -492001
rect -50 -492143 -34 -492109
rect 34 -492143 50 -492109
rect -96 -492193 -62 -492177
rect -96 -493185 -62 -493169
rect 62 -492193 96 -492177
rect 62 -493185 96 -493169
rect -50 -493253 -34 -493219
rect 34 -493253 50 -493219
rect -50 -493361 -34 -493327
rect 34 -493361 50 -493327
rect -96 -493411 -62 -493395
rect -96 -494403 -62 -494387
rect 62 -493411 96 -493395
rect 62 -494403 96 -494387
rect -50 -494471 -34 -494437
rect 34 -494471 50 -494437
rect -50 -494579 -34 -494545
rect 34 -494579 50 -494545
rect -96 -494629 -62 -494613
rect -96 -495621 -62 -495605
rect 62 -494629 96 -494613
rect 62 -495621 96 -495605
rect -50 -495689 -34 -495655
rect 34 -495689 50 -495655
rect -50 -495797 -34 -495763
rect 34 -495797 50 -495763
rect -96 -495847 -62 -495831
rect -96 -496839 -62 -496823
rect 62 -495847 96 -495831
rect 62 -496839 96 -496823
rect -50 -496907 -34 -496873
rect 34 -496907 50 -496873
rect -50 -497015 -34 -496981
rect 34 -497015 50 -496981
rect -96 -497065 -62 -497049
rect -96 -498057 -62 -498041
rect 62 -497065 96 -497049
rect 62 -498057 96 -498041
rect -50 -498125 -34 -498091
rect 34 -498125 50 -498091
rect -50 -498233 -34 -498199
rect 34 -498233 50 -498199
rect -96 -498283 -62 -498267
rect -96 -499275 -62 -499259
rect 62 -498283 96 -498267
rect 62 -499275 96 -499259
rect -50 -499343 -34 -499309
rect 34 -499343 50 -499309
rect -50 -499451 -34 -499417
rect 34 -499451 50 -499417
rect -96 -499501 -62 -499485
rect -96 -500493 -62 -500477
rect 62 -499501 96 -499485
rect 62 -500493 96 -500477
rect -50 -500561 -34 -500527
rect 34 -500561 50 -500527
rect -50 -500669 -34 -500635
rect 34 -500669 50 -500635
rect -96 -500719 -62 -500703
rect -96 -501711 -62 -501695
rect 62 -500719 96 -500703
rect 62 -501711 96 -501695
rect -50 -501779 -34 -501745
rect 34 -501779 50 -501745
rect -50 -501887 -34 -501853
rect 34 -501887 50 -501853
rect -96 -501937 -62 -501921
rect -96 -502929 -62 -502913
rect 62 -501937 96 -501921
rect 62 -502929 96 -502913
rect -50 -502997 -34 -502963
rect 34 -502997 50 -502963
rect -50 -503105 -34 -503071
rect 34 -503105 50 -503071
rect -96 -503155 -62 -503139
rect -96 -504147 -62 -504131
rect 62 -503155 96 -503139
rect 62 -504147 96 -504131
rect -50 -504215 -34 -504181
rect 34 -504215 50 -504181
rect -50 -504323 -34 -504289
rect 34 -504323 50 -504289
rect -96 -504373 -62 -504357
rect -96 -505365 -62 -505349
rect 62 -504373 96 -504357
rect 62 -505365 96 -505349
rect -50 -505433 -34 -505399
rect 34 -505433 50 -505399
rect -50 -505541 -34 -505507
rect 34 -505541 50 -505507
rect -96 -505591 -62 -505575
rect -96 -506583 -62 -506567
rect 62 -505591 96 -505575
rect 62 -506583 96 -506567
rect -50 -506651 -34 -506617
rect 34 -506651 50 -506617
rect -50 -506759 -34 -506725
rect 34 -506759 50 -506725
rect -96 -506809 -62 -506793
rect -96 -507801 -62 -507785
rect 62 -506809 96 -506793
rect 62 -507801 96 -507785
rect -50 -507869 -34 -507835
rect 34 -507869 50 -507835
rect -50 -507977 -34 -507943
rect 34 -507977 50 -507943
rect -96 -508027 -62 -508011
rect -96 -509019 -62 -509003
rect 62 -508027 96 -508011
rect 62 -509019 96 -509003
rect -50 -509087 -34 -509053
rect 34 -509087 50 -509053
rect -50 -509195 -34 -509161
rect 34 -509195 50 -509161
rect -96 -509245 -62 -509229
rect -96 -510237 -62 -510221
rect 62 -509245 96 -509229
rect 62 -510237 96 -510221
rect -50 -510305 -34 -510271
rect 34 -510305 50 -510271
rect -50 -510413 -34 -510379
rect 34 -510413 50 -510379
rect -96 -510463 -62 -510447
rect -96 -511455 -62 -511439
rect 62 -510463 96 -510447
rect 62 -511455 96 -511439
rect -50 -511523 -34 -511489
rect 34 -511523 50 -511489
rect -50 -511631 -34 -511597
rect 34 -511631 50 -511597
rect -96 -511681 -62 -511665
rect -96 -512673 -62 -512657
rect 62 -511681 96 -511665
rect 62 -512673 96 -512657
rect -50 -512741 -34 -512707
rect 34 -512741 50 -512707
rect -50 -512849 -34 -512815
rect 34 -512849 50 -512815
rect -96 -512899 -62 -512883
rect -96 -513891 -62 -513875
rect 62 -512899 96 -512883
rect 62 -513891 96 -513875
rect -50 -513959 -34 -513925
rect 34 -513959 50 -513925
rect -50 -514067 -34 -514033
rect 34 -514067 50 -514033
rect -96 -514117 -62 -514101
rect -96 -515109 -62 -515093
rect 62 -514117 96 -514101
rect 62 -515109 96 -515093
rect -50 -515177 -34 -515143
rect 34 -515177 50 -515143
rect -50 -515285 -34 -515251
rect 34 -515285 50 -515251
rect -96 -515335 -62 -515319
rect -96 -516327 -62 -516311
rect 62 -515335 96 -515319
rect 62 -516327 96 -516311
rect -50 -516395 -34 -516361
rect 34 -516395 50 -516361
rect -50 -516503 -34 -516469
rect 34 -516503 50 -516469
rect -96 -516553 -62 -516537
rect -96 -517545 -62 -517529
rect 62 -516553 96 -516537
rect 62 -517545 96 -517529
rect -50 -517613 -34 -517579
rect 34 -517613 50 -517579
rect -50 -517721 -34 -517687
rect 34 -517721 50 -517687
rect -96 -517771 -62 -517755
rect -96 -518763 -62 -518747
rect 62 -517771 96 -517755
rect 62 -518763 96 -518747
rect -50 -518831 -34 -518797
rect 34 -518831 50 -518797
rect -50 -518939 -34 -518905
rect 34 -518939 50 -518905
rect -96 -518989 -62 -518973
rect -96 -519981 -62 -519965
rect 62 -518989 96 -518973
rect 62 -519981 96 -519965
rect -50 -520049 -34 -520015
rect 34 -520049 50 -520015
rect -50 -520157 -34 -520123
rect 34 -520157 50 -520123
rect -96 -520207 -62 -520191
rect -96 -521199 -62 -521183
rect 62 -520207 96 -520191
rect 62 -521199 96 -521183
rect -50 -521267 -34 -521233
rect 34 -521267 50 -521233
rect -50 -521375 -34 -521341
rect 34 -521375 50 -521341
rect -96 -521425 -62 -521409
rect -96 -522417 -62 -522401
rect 62 -521425 96 -521409
rect 62 -522417 96 -522401
rect -50 -522485 -34 -522451
rect 34 -522485 50 -522451
rect -50 -522593 -34 -522559
rect 34 -522593 50 -522559
rect -96 -522643 -62 -522627
rect -96 -523635 -62 -523619
rect 62 -522643 96 -522627
rect 62 -523635 96 -523619
rect -50 -523703 -34 -523669
rect 34 -523703 50 -523669
rect -50 -523811 -34 -523777
rect 34 -523811 50 -523777
rect -96 -523861 -62 -523845
rect -96 -524853 -62 -524837
rect 62 -523861 96 -523845
rect 62 -524853 96 -524837
rect -50 -524921 -34 -524887
rect 34 -524921 50 -524887
rect -50 -525029 -34 -524995
rect 34 -525029 50 -524995
rect -96 -525079 -62 -525063
rect -96 -526071 -62 -526055
rect 62 -525079 96 -525063
rect 62 -526071 96 -526055
rect -50 -526139 -34 -526105
rect 34 -526139 50 -526105
rect -50 -526247 -34 -526213
rect 34 -526247 50 -526213
rect -96 -526297 -62 -526281
rect -96 -527289 -62 -527273
rect 62 -526297 96 -526281
rect 62 -527289 96 -527273
rect -50 -527357 -34 -527323
rect 34 -527357 50 -527323
rect -50 -527465 -34 -527431
rect 34 -527465 50 -527431
rect -96 -527515 -62 -527499
rect -96 -528507 -62 -528491
rect 62 -527515 96 -527499
rect 62 -528507 96 -528491
rect -50 -528575 -34 -528541
rect 34 -528575 50 -528541
rect -50 -528683 -34 -528649
rect 34 -528683 50 -528649
rect -96 -528733 -62 -528717
rect -96 -529725 -62 -529709
rect 62 -528733 96 -528717
rect 62 -529725 96 -529709
rect -50 -529793 -34 -529759
rect 34 -529793 50 -529759
rect -50 -529901 -34 -529867
rect 34 -529901 50 -529867
rect -96 -529951 -62 -529935
rect -96 -530943 -62 -530927
rect 62 -529951 96 -529935
rect 62 -530943 96 -530927
rect -50 -531011 -34 -530977
rect 34 -531011 50 -530977
rect -50 -531119 -34 -531085
rect 34 -531119 50 -531085
rect -96 -531169 -62 -531153
rect -96 -532161 -62 -532145
rect 62 -531169 96 -531153
rect 62 -532161 96 -532145
rect -50 -532229 -34 -532195
rect 34 -532229 50 -532195
rect -50 -532337 -34 -532303
rect 34 -532337 50 -532303
rect -96 -532387 -62 -532371
rect -96 -533379 -62 -533363
rect 62 -532387 96 -532371
rect 62 -533379 96 -533363
rect -50 -533447 -34 -533413
rect 34 -533447 50 -533413
rect -50 -533555 -34 -533521
rect 34 -533555 50 -533521
rect -96 -533605 -62 -533589
rect -96 -534597 -62 -534581
rect 62 -533605 96 -533589
rect 62 -534597 96 -534581
rect -50 -534665 -34 -534631
rect 34 -534665 50 -534631
rect -50 -534773 -34 -534739
rect 34 -534773 50 -534739
rect -96 -534823 -62 -534807
rect -96 -535815 -62 -535799
rect 62 -534823 96 -534807
rect 62 -535815 96 -535799
rect -50 -535883 -34 -535849
rect 34 -535883 50 -535849
rect -50 -535991 -34 -535957
rect 34 -535991 50 -535957
rect -96 -536041 -62 -536025
rect -96 -537033 -62 -537017
rect 62 -536041 96 -536025
rect 62 -537033 96 -537017
rect -50 -537101 -34 -537067
rect 34 -537101 50 -537067
rect -50 -537209 -34 -537175
rect 34 -537209 50 -537175
rect -96 -537259 -62 -537243
rect -96 -538251 -62 -538235
rect 62 -537259 96 -537243
rect 62 -538251 96 -538235
rect -50 -538319 -34 -538285
rect 34 -538319 50 -538285
rect -50 -538427 -34 -538393
rect 34 -538427 50 -538393
rect -96 -538477 -62 -538461
rect -96 -539469 -62 -539453
rect 62 -538477 96 -538461
rect 62 -539469 96 -539453
rect -50 -539537 -34 -539503
rect 34 -539537 50 -539503
rect -50 -539645 -34 -539611
rect 34 -539645 50 -539611
rect -96 -539695 -62 -539679
rect -96 -540687 -62 -540671
rect 62 -539695 96 -539679
rect 62 -540687 96 -540671
rect -50 -540755 -34 -540721
rect 34 -540755 50 -540721
rect -50 -540863 -34 -540829
rect 34 -540863 50 -540829
rect -96 -540913 -62 -540897
rect -96 -541905 -62 -541889
rect 62 -540913 96 -540897
rect 62 -541905 96 -541889
rect -50 -541973 -34 -541939
rect 34 -541973 50 -541939
rect -50 -542081 -34 -542047
rect 34 -542081 50 -542047
rect -96 -542131 -62 -542115
rect -96 -543123 -62 -543107
rect 62 -542131 96 -542115
rect 62 -543123 96 -543107
rect -50 -543191 -34 -543157
rect 34 -543191 50 -543157
rect -50 -543299 -34 -543265
rect 34 -543299 50 -543265
rect -96 -543349 -62 -543333
rect -96 -544341 -62 -544325
rect 62 -543349 96 -543333
rect 62 -544341 96 -544325
rect -50 -544409 -34 -544375
rect 34 -544409 50 -544375
rect -50 -544517 -34 -544483
rect 34 -544517 50 -544483
rect -96 -544567 -62 -544551
rect -96 -545559 -62 -545543
rect 62 -544567 96 -544551
rect 62 -545559 96 -545543
rect -50 -545627 -34 -545593
rect 34 -545627 50 -545593
rect -50 -545735 -34 -545701
rect 34 -545735 50 -545701
rect -96 -545785 -62 -545769
rect -96 -546777 -62 -546761
rect 62 -545785 96 -545769
rect 62 -546777 96 -546761
rect -50 -546845 -34 -546811
rect 34 -546845 50 -546811
rect -50 -546953 -34 -546919
rect 34 -546953 50 -546919
rect -96 -547003 -62 -546987
rect -96 -547995 -62 -547979
rect 62 -547003 96 -546987
rect 62 -547995 96 -547979
rect -50 -548063 -34 -548029
rect 34 -548063 50 -548029
rect -50 -548171 -34 -548137
rect 34 -548171 50 -548137
rect -96 -548221 -62 -548205
rect -96 -549213 -62 -549197
rect 62 -548221 96 -548205
rect 62 -549213 96 -549197
rect -50 -549281 -34 -549247
rect 34 -549281 50 -549247
rect -50 -549389 -34 -549355
rect 34 -549389 50 -549355
rect -96 -549439 -62 -549423
rect -96 -550431 -62 -550415
rect 62 -549439 96 -549423
rect 62 -550431 96 -550415
rect -50 -550499 -34 -550465
rect 34 -550499 50 -550465
rect -50 -550607 -34 -550573
rect 34 -550607 50 -550573
rect -96 -550657 -62 -550641
rect -96 -551649 -62 -551633
rect 62 -550657 96 -550641
rect 62 -551649 96 -551633
rect -50 -551717 -34 -551683
rect 34 -551717 50 -551683
rect -50 -551825 -34 -551791
rect 34 -551825 50 -551791
rect -96 -551875 -62 -551859
rect -96 -552867 -62 -552851
rect 62 -551875 96 -551859
rect 62 -552867 96 -552851
rect -50 -552935 -34 -552901
rect 34 -552935 50 -552901
rect -50 -553043 -34 -553009
rect 34 -553043 50 -553009
rect -96 -553093 -62 -553077
rect -96 -554085 -62 -554069
rect 62 -553093 96 -553077
rect 62 -554085 96 -554069
rect -50 -554153 -34 -554119
rect 34 -554153 50 -554119
rect -50 -554261 -34 -554227
rect 34 -554261 50 -554227
rect -96 -554311 -62 -554295
rect -96 -555303 -62 -555287
rect 62 -554311 96 -554295
rect 62 -555303 96 -555287
rect -50 -555371 -34 -555337
rect 34 -555371 50 -555337
rect -50 -555479 -34 -555445
rect 34 -555479 50 -555445
rect -96 -555529 -62 -555513
rect -96 -556521 -62 -556505
rect 62 -555529 96 -555513
rect 62 -556521 96 -556505
rect -50 -556589 -34 -556555
rect 34 -556589 50 -556555
rect -50 -556697 -34 -556663
rect 34 -556697 50 -556663
rect -96 -556747 -62 -556731
rect -96 -557739 -62 -557723
rect 62 -556747 96 -556731
rect 62 -557739 96 -557723
rect -50 -557807 -34 -557773
rect 34 -557807 50 -557773
rect -50 -557915 -34 -557881
rect 34 -557915 50 -557881
rect -96 -557965 -62 -557949
rect -96 -558957 -62 -558941
rect 62 -557965 96 -557949
rect 62 -558957 96 -558941
rect -50 -559025 -34 -558991
rect 34 -559025 50 -558991
rect -50 -559133 -34 -559099
rect 34 -559133 50 -559099
rect -96 -559183 -62 -559167
rect -96 -560175 -62 -560159
rect 62 -559183 96 -559167
rect 62 -560175 96 -560159
rect -50 -560243 -34 -560209
rect 34 -560243 50 -560209
rect -50 -560351 -34 -560317
rect 34 -560351 50 -560317
rect -96 -560401 -62 -560385
rect -96 -561393 -62 -561377
rect 62 -560401 96 -560385
rect 62 -561393 96 -561377
rect -50 -561461 -34 -561427
rect 34 -561461 50 -561427
rect -50 -561569 -34 -561535
rect 34 -561569 50 -561535
rect -96 -561619 -62 -561603
rect -96 -562611 -62 -562595
rect 62 -561619 96 -561603
rect 62 -562611 96 -562595
rect -50 -562679 -34 -562645
rect 34 -562679 50 -562645
rect -50 -562787 -34 -562753
rect 34 -562787 50 -562753
rect -96 -562837 -62 -562821
rect -96 -563829 -62 -563813
rect 62 -562837 96 -562821
rect 62 -563829 96 -563813
rect -50 -563897 -34 -563863
rect 34 -563897 50 -563863
rect -50 -564005 -34 -563971
rect 34 -564005 50 -563971
rect -96 -564055 -62 -564039
rect -96 -565047 -62 -565031
rect 62 -564055 96 -564039
rect 62 -565047 96 -565031
rect -50 -565115 -34 -565081
rect 34 -565115 50 -565081
rect -50 -565223 -34 -565189
rect 34 -565223 50 -565189
rect -96 -565273 -62 -565257
rect -96 -566265 -62 -566249
rect 62 -565273 96 -565257
rect 62 -566265 96 -566249
rect -50 -566333 -34 -566299
rect 34 -566333 50 -566299
rect -50 -566441 -34 -566407
rect 34 -566441 50 -566407
rect -96 -566491 -62 -566475
rect -96 -567483 -62 -567467
rect 62 -566491 96 -566475
rect 62 -567483 96 -567467
rect -50 -567551 -34 -567517
rect 34 -567551 50 -567517
rect -50 -567659 -34 -567625
rect 34 -567659 50 -567625
rect -96 -567709 -62 -567693
rect -96 -568701 -62 -568685
rect 62 -567709 96 -567693
rect 62 -568701 96 -568685
rect -50 -568769 -34 -568735
rect 34 -568769 50 -568735
rect -50 -568877 -34 -568843
rect 34 -568877 50 -568843
rect -96 -568927 -62 -568911
rect -96 -569919 -62 -569903
rect 62 -568927 96 -568911
rect 62 -569919 96 -569903
rect -50 -569987 -34 -569953
rect 34 -569987 50 -569953
rect -50 -570095 -34 -570061
rect 34 -570095 50 -570061
rect -96 -570145 -62 -570129
rect -96 -571137 -62 -571121
rect 62 -570145 96 -570129
rect 62 -571137 96 -571121
rect -50 -571205 -34 -571171
rect 34 -571205 50 -571171
rect -50 -571313 -34 -571279
rect 34 -571313 50 -571279
rect -96 -571363 -62 -571347
rect -96 -572355 -62 -572339
rect 62 -571363 96 -571347
rect 62 -572355 96 -572339
rect -50 -572423 -34 -572389
rect 34 -572423 50 -572389
rect -50 -572531 -34 -572497
rect 34 -572531 50 -572497
rect -96 -572581 -62 -572565
rect -96 -573573 -62 -573557
rect 62 -572581 96 -572565
rect 62 -573573 96 -573557
rect -50 -573641 -34 -573607
rect 34 -573641 50 -573607
rect -50 -573749 -34 -573715
rect 34 -573749 50 -573715
rect -96 -573799 -62 -573783
rect -96 -574791 -62 -574775
rect 62 -573799 96 -573783
rect 62 -574791 96 -574775
rect -50 -574859 -34 -574825
rect 34 -574859 50 -574825
rect -50 -574967 -34 -574933
rect 34 -574967 50 -574933
rect -96 -575017 -62 -575001
rect -96 -576009 -62 -575993
rect 62 -575017 96 -575001
rect 62 -576009 96 -575993
rect -50 -576077 -34 -576043
rect 34 -576077 50 -576043
rect -50 -576185 -34 -576151
rect 34 -576185 50 -576151
rect -96 -576235 -62 -576219
rect -96 -577227 -62 -577211
rect 62 -576235 96 -576219
rect 62 -577227 96 -577211
rect -50 -577295 -34 -577261
rect 34 -577295 50 -577261
rect -50 -577403 -34 -577369
rect 34 -577403 50 -577369
rect -96 -577453 -62 -577437
rect -96 -578445 -62 -578429
rect 62 -577453 96 -577437
rect 62 -578445 96 -578429
rect -50 -578513 -34 -578479
rect 34 -578513 50 -578479
rect -50 -578621 -34 -578587
rect 34 -578621 50 -578587
rect -96 -578671 -62 -578655
rect -96 -579663 -62 -579647
rect 62 -578671 96 -578655
rect 62 -579663 96 -579647
rect -50 -579731 -34 -579697
rect 34 -579731 50 -579697
rect -50 -579839 -34 -579805
rect 34 -579839 50 -579805
rect -96 -579889 -62 -579873
rect -96 -580881 -62 -580865
rect 62 -579889 96 -579873
rect 62 -580881 96 -580865
rect -50 -580949 -34 -580915
rect 34 -580949 50 -580915
rect -50 -581057 -34 -581023
rect 34 -581057 50 -581023
rect -96 -581107 -62 -581091
rect -96 -582099 -62 -582083
rect 62 -581107 96 -581091
rect 62 -582099 96 -582083
rect -50 -582167 -34 -582133
rect 34 -582167 50 -582133
rect -50 -582275 -34 -582241
rect 34 -582275 50 -582241
rect -96 -582325 -62 -582309
rect -96 -583317 -62 -583301
rect 62 -582325 96 -582309
rect 62 -583317 96 -583301
rect -50 -583385 -34 -583351
rect 34 -583385 50 -583351
rect -50 -583493 -34 -583459
rect 34 -583493 50 -583459
rect -96 -583543 -62 -583527
rect -96 -584535 -62 -584519
rect 62 -583543 96 -583527
rect 62 -584535 96 -584519
rect -50 -584603 -34 -584569
rect 34 -584603 50 -584569
rect -50 -584711 -34 -584677
rect 34 -584711 50 -584677
rect -96 -584761 -62 -584745
rect -96 -585753 -62 -585737
rect 62 -584761 96 -584745
rect 62 -585753 96 -585737
rect -50 -585821 -34 -585787
rect 34 -585821 50 -585787
rect -50 -585929 -34 -585895
rect 34 -585929 50 -585895
rect -96 -585979 -62 -585963
rect -96 -586971 -62 -586955
rect 62 -585979 96 -585963
rect 62 -586971 96 -586955
rect -50 -587039 -34 -587005
rect 34 -587039 50 -587005
rect -50 -587147 -34 -587113
rect 34 -587147 50 -587113
rect -96 -587197 -62 -587181
rect -96 -588189 -62 -588173
rect 62 -587197 96 -587181
rect 62 -588189 96 -588173
rect -50 -588257 -34 -588223
rect 34 -588257 50 -588223
rect -50 -588365 -34 -588331
rect 34 -588365 50 -588331
rect -96 -588415 -62 -588399
rect -96 -589407 -62 -589391
rect 62 -588415 96 -588399
rect 62 -589407 96 -589391
rect -50 -589475 -34 -589441
rect 34 -589475 50 -589441
rect -50 -589583 -34 -589549
rect 34 -589583 50 -589549
rect -96 -589633 -62 -589617
rect -96 -590625 -62 -590609
rect 62 -589633 96 -589617
rect 62 -590625 96 -590609
rect -50 -590693 -34 -590659
rect 34 -590693 50 -590659
rect -50 -590801 -34 -590767
rect 34 -590801 50 -590767
rect -96 -590851 -62 -590835
rect -96 -591843 -62 -591827
rect 62 -590851 96 -590835
rect 62 -591843 96 -591827
rect -50 -591911 -34 -591877
rect 34 -591911 50 -591877
rect -50 -592019 -34 -591985
rect 34 -592019 50 -591985
rect -96 -592069 -62 -592053
rect -96 -593061 -62 -593045
rect 62 -592069 96 -592053
rect 62 -593061 96 -593045
rect -50 -593129 -34 -593095
rect 34 -593129 50 -593095
rect -50 -593237 -34 -593203
rect 34 -593237 50 -593203
rect -96 -593287 -62 -593271
rect -96 -594279 -62 -594263
rect 62 -593287 96 -593271
rect 62 -594279 96 -594263
rect -50 -594347 -34 -594313
rect 34 -594347 50 -594313
rect -50 -594455 -34 -594421
rect 34 -594455 50 -594421
rect -96 -594505 -62 -594489
rect -96 -595497 -62 -595481
rect 62 -594505 96 -594489
rect 62 -595497 96 -595481
rect -50 -595565 -34 -595531
rect 34 -595565 50 -595531
rect -50 -595673 -34 -595639
rect 34 -595673 50 -595639
rect -96 -595723 -62 -595707
rect -96 -596715 -62 -596699
rect 62 -595723 96 -595707
rect 62 -596715 96 -596699
rect -50 -596783 -34 -596749
rect 34 -596783 50 -596749
rect -50 -596891 -34 -596857
rect 34 -596891 50 -596857
rect -96 -596941 -62 -596925
rect -96 -597933 -62 -597917
rect 62 -596941 96 -596925
rect 62 -597933 96 -597917
rect -50 -598001 -34 -597967
rect 34 -598001 50 -597967
rect -50 -598109 -34 -598075
rect 34 -598109 50 -598075
rect -96 -598159 -62 -598143
rect -96 -599151 -62 -599135
rect 62 -598159 96 -598143
rect 62 -599151 96 -599135
rect -50 -599219 -34 -599185
rect 34 -599219 50 -599185
rect -50 -599327 -34 -599293
rect 34 -599327 50 -599293
rect -96 -599377 -62 -599361
rect -96 -600369 -62 -600353
rect 62 -599377 96 -599361
rect 62 -600369 96 -600353
rect -50 -600437 -34 -600403
rect 34 -600437 50 -600403
rect -50 -600545 -34 -600511
rect 34 -600545 50 -600511
rect -96 -600595 -62 -600579
rect -96 -601587 -62 -601571
rect 62 -600595 96 -600579
rect 62 -601587 96 -601571
rect -50 -601655 -34 -601621
rect 34 -601655 50 -601621
rect -50 -601763 -34 -601729
rect 34 -601763 50 -601729
rect -96 -601813 -62 -601797
rect -96 -602805 -62 -602789
rect 62 -601813 96 -601797
rect 62 -602805 96 -602789
rect -50 -602873 -34 -602839
rect 34 -602873 50 -602839
rect -50 -602981 -34 -602947
rect 34 -602981 50 -602947
rect -96 -603031 -62 -603015
rect -96 -604023 -62 -604007
rect 62 -603031 96 -603015
rect 62 -604023 96 -604007
rect -50 -604091 -34 -604057
rect 34 -604091 50 -604057
rect -50 -604199 -34 -604165
rect 34 -604199 50 -604165
rect -96 -604249 -62 -604233
rect -96 -605241 -62 -605225
rect 62 -604249 96 -604233
rect 62 -605241 96 -605225
rect -50 -605309 -34 -605275
rect 34 -605309 50 -605275
rect -50 -605417 -34 -605383
rect 34 -605417 50 -605383
rect -96 -605467 -62 -605451
rect -96 -606459 -62 -606443
rect 62 -605467 96 -605451
rect 62 -606459 96 -606443
rect -50 -606527 -34 -606493
rect 34 -606527 50 -606493
rect -50 -606635 -34 -606601
rect 34 -606635 50 -606601
rect -96 -606685 -62 -606669
rect -96 -607677 -62 -607661
rect 62 -606685 96 -606669
rect 62 -607677 96 -607661
rect -50 -607745 -34 -607711
rect 34 -607745 50 -607711
rect -50 -607853 -34 -607819
rect 34 -607853 50 -607819
rect -96 -607903 -62 -607887
rect -96 -608895 -62 -608879
rect 62 -607903 96 -607887
rect 62 -608895 96 -608879
rect -50 -608963 -34 -608929
rect 34 -608963 50 -608929
rect -230 -609067 -196 -609005
rect 196 -609067 230 -609005
rect -230 -609101 -134 -609067
rect 134 -609101 230 -609067
<< viali >>
rect -34 608929 34 608963
rect -96 607903 -62 608879
rect 62 607903 96 608879
rect -34 607819 34 607853
rect -34 607711 34 607745
rect -96 606685 -62 607661
rect 62 606685 96 607661
rect -34 606601 34 606635
rect -34 606493 34 606527
rect -96 605467 -62 606443
rect 62 605467 96 606443
rect -34 605383 34 605417
rect -34 605275 34 605309
rect -96 604249 -62 605225
rect 62 604249 96 605225
rect -34 604165 34 604199
rect -34 604057 34 604091
rect -96 603031 -62 604007
rect 62 603031 96 604007
rect -34 602947 34 602981
rect -34 602839 34 602873
rect -96 601813 -62 602789
rect 62 601813 96 602789
rect -34 601729 34 601763
rect -34 601621 34 601655
rect -96 600595 -62 601571
rect 62 600595 96 601571
rect -34 600511 34 600545
rect -34 600403 34 600437
rect -96 599377 -62 600353
rect 62 599377 96 600353
rect -34 599293 34 599327
rect -34 599185 34 599219
rect -96 598159 -62 599135
rect 62 598159 96 599135
rect -34 598075 34 598109
rect -34 597967 34 598001
rect -96 596941 -62 597917
rect 62 596941 96 597917
rect -34 596857 34 596891
rect -34 596749 34 596783
rect -96 595723 -62 596699
rect 62 595723 96 596699
rect -34 595639 34 595673
rect -34 595531 34 595565
rect -96 594505 -62 595481
rect 62 594505 96 595481
rect -34 594421 34 594455
rect -34 594313 34 594347
rect -96 593287 -62 594263
rect 62 593287 96 594263
rect -34 593203 34 593237
rect -34 593095 34 593129
rect -96 592069 -62 593045
rect 62 592069 96 593045
rect -34 591985 34 592019
rect -34 591877 34 591911
rect -96 590851 -62 591827
rect 62 590851 96 591827
rect -34 590767 34 590801
rect -34 590659 34 590693
rect -96 589633 -62 590609
rect 62 589633 96 590609
rect -34 589549 34 589583
rect -34 589441 34 589475
rect -96 588415 -62 589391
rect 62 588415 96 589391
rect -34 588331 34 588365
rect -34 588223 34 588257
rect -96 587197 -62 588173
rect 62 587197 96 588173
rect -34 587113 34 587147
rect -34 587005 34 587039
rect -96 585979 -62 586955
rect 62 585979 96 586955
rect -34 585895 34 585929
rect -34 585787 34 585821
rect -96 584761 -62 585737
rect 62 584761 96 585737
rect -34 584677 34 584711
rect -34 584569 34 584603
rect -96 583543 -62 584519
rect 62 583543 96 584519
rect -34 583459 34 583493
rect -34 583351 34 583385
rect -96 582325 -62 583301
rect 62 582325 96 583301
rect -34 582241 34 582275
rect -34 582133 34 582167
rect -96 581107 -62 582083
rect 62 581107 96 582083
rect -34 581023 34 581057
rect -34 580915 34 580949
rect -96 579889 -62 580865
rect 62 579889 96 580865
rect -34 579805 34 579839
rect -34 579697 34 579731
rect -96 578671 -62 579647
rect 62 578671 96 579647
rect -34 578587 34 578621
rect -34 578479 34 578513
rect -96 577453 -62 578429
rect 62 577453 96 578429
rect -34 577369 34 577403
rect -34 577261 34 577295
rect -96 576235 -62 577211
rect 62 576235 96 577211
rect -34 576151 34 576185
rect -34 576043 34 576077
rect -96 575017 -62 575993
rect 62 575017 96 575993
rect -34 574933 34 574967
rect -34 574825 34 574859
rect -96 573799 -62 574775
rect 62 573799 96 574775
rect -34 573715 34 573749
rect -34 573607 34 573641
rect -96 572581 -62 573557
rect 62 572581 96 573557
rect -34 572497 34 572531
rect -34 572389 34 572423
rect -96 571363 -62 572339
rect 62 571363 96 572339
rect -34 571279 34 571313
rect -34 571171 34 571205
rect -96 570145 -62 571121
rect 62 570145 96 571121
rect -34 570061 34 570095
rect -34 569953 34 569987
rect -96 568927 -62 569903
rect 62 568927 96 569903
rect -34 568843 34 568877
rect -34 568735 34 568769
rect -96 567709 -62 568685
rect 62 567709 96 568685
rect -34 567625 34 567659
rect -34 567517 34 567551
rect -96 566491 -62 567467
rect 62 566491 96 567467
rect -34 566407 34 566441
rect -34 566299 34 566333
rect -96 565273 -62 566249
rect 62 565273 96 566249
rect -34 565189 34 565223
rect -34 565081 34 565115
rect -96 564055 -62 565031
rect 62 564055 96 565031
rect -34 563971 34 564005
rect -34 563863 34 563897
rect -96 562837 -62 563813
rect 62 562837 96 563813
rect -34 562753 34 562787
rect -34 562645 34 562679
rect -96 561619 -62 562595
rect 62 561619 96 562595
rect -34 561535 34 561569
rect -34 561427 34 561461
rect -96 560401 -62 561377
rect 62 560401 96 561377
rect -34 560317 34 560351
rect -34 560209 34 560243
rect -96 559183 -62 560159
rect 62 559183 96 560159
rect -34 559099 34 559133
rect -34 558991 34 559025
rect -96 557965 -62 558941
rect 62 557965 96 558941
rect -34 557881 34 557915
rect -34 557773 34 557807
rect -96 556747 -62 557723
rect 62 556747 96 557723
rect -34 556663 34 556697
rect -34 556555 34 556589
rect -96 555529 -62 556505
rect 62 555529 96 556505
rect -34 555445 34 555479
rect -34 555337 34 555371
rect -96 554311 -62 555287
rect 62 554311 96 555287
rect -34 554227 34 554261
rect -34 554119 34 554153
rect -96 553093 -62 554069
rect 62 553093 96 554069
rect -34 553009 34 553043
rect -34 552901 34 552935
rect -96 551875 -62 552851
rect 62 551875 96 552851
rect -34 551791 34 551825
rect -34 551683 34 551717
rect -96 550657 -62 551633
rect 62 550657 96 551633
rect -34 550573 34 550607
rect -34 550465 34 550499
rect -96 549439 -62 550415
rect 62 549439 96 550415
rect -34 549355 34 549389
rect -34 549247 34 549281
rect -96 548221 -62 549197
rect 62 548221 96 549197
rect -34 548137 34 548171
rect -34 548029 34 548063
rect -96 547003 -62 547979
rect 62 547003 96 547979
rect -34 546919 34 546953
rect -34 546811 34 546845
rect -96 545785 -62 546761
rect 62 545785 96 546761
rect -34 545701 34 545735
rect -34 545593 34 545627
rect -96 544567 -62 545543
rect 62 544567 96 545543
rect -34 544483 34 544517
rect -34 544375 34 544409
rect -96 543349 -62 544325
rect 62 543349 96 544325
rect -34 543265 34 543299
rect -34 543157 34 543191
rect -96 542131 -62 543107
rect 62 542131 96 543107
rect -34 542047 34 542081
rect -34 541939 34 541973
rect -96 540913 -62 541889
rect 62 540913 96 541889
rect -34 540829 34 540863
rect -34 540721 34 540755
rect -96 539695 -62 540671
rect 62 539695 96 540671
rect -34 539611 34 539645
rect -34 539503 34 539537
rect -96 538477 -62 539453
rect 62 538477 96 539453
rect -34 538393 34 538427
rect -34 538285 34 538319
rect -96 537259 -62 538235
rect 62 537259 96 538235
rect -34 537175 34 537209
rect -34 537067 34 537101
rect -96 536041 -62 537017
rect 62 536041 96 537017
rect -34 535957 34 535991
rect -34 535849 34 535883
rect -96 534823 -62 535799
rect 62 534823 96 535799
rect -34 534739 34 534773
rect -34 534631 34 534665
rect -96 533605 -62 534581
rect 62 533605 96 534581
rect -34 533521 34 533555
rect -34 533413 34 533447
rect -96 532387 -62 533363
rect 62 532387 96 533363
rect -34 532303 34 532337
rect -34 532195 34 532229
rect -96 531169 -62 532145
rect 62 531169 96 532145
rect -34 531085 34 531119
rect -34 530977 34 531011
rect -96 529951 -62 530927
rect 62 529951 96 530927
rect -34 529867 34 529901
rect -34 529759 34 529793
rect -96 528733 -62 529709
rect 62 528733 96 529709
rect -34 528649 34 528683
rect -34 528541 34 528575
rect -96 527515 -62 528491
rect 62 527515 96 528491
rect -34 527431 34 527465
rect -34 527323 34 527357
rect -96 526297 -62 527273
rect 62 526297 96 527273
rect -34 526213 34 526247
rect -34 526105 34 526139
rect -96 525079 -62 526055
rect 62 525079 96 526055
rect -34 524995 34 525029
rect -34 524887 34 524921
rect -96 523861 -62 524837
rect 62 523861 96 524837
rect -34 523777 34 523811
rect -34 523669 34 523703
rect -96 522643 -62 523619
rect 62 522643 96 523619
rect -34 522559 34 522593
rect -34 522451 34 522485
rect -96 521425 -62 522401
rect 62 521425 96 522401
rect -34 521341 34 521375
rect -34 521233 34 521267
rect -96 520207 -62 521183
rect 62 520207 96 521183
rect -34 520123 34 520157
rect -34 520015 34 520049
rect -96 518989 -62 519965
rect 62 518989 96 519965
rect -34 518905 34 518939
rect -34 518797 34 518831
rect -96 517771 -62 518747
rect 62 517771 96 518747
rect -34 517687 34 517721
rect -34 517579 34 517613
rect -96 516553 -62 517529
rect 62 516553 96 517529
rect -34 516469 34 516503
rect -34 516361 34 516395
rect -96 515335 -62 516311
rect 62 515335 96 516311
rect -34 515251 34 515285
rect -34 515143 34 515177
rect -96 514117 -62 515093
rect 62 514117 96 515093
rect -34 514033 34 514067
rect -34 513925 34 513959
rect -96 512899 -62 513875
rect 62 512899 96 513875
rect -34 512815 34 512849
rect -34 512707 34 512741
rect -96 511681 -62 512657
rect 62 511681 96 512657
rect -34 511597 34 511631
rect -34 511489 34 511523
rect -96 510463 -62 511439
rect 62 510463 96 511439
rect -34 510379 34 510413
rect -34 510271 34 510305
rect -96 509245 -62 510221
rect 62 509245 96 510221
rect -34 509161 34 509195
rect -34 509053 34 509087
rect -96 508027 -62 509003
rect 62 508027 96 509003
rect -34 507943 34 507977
rect -34 507835 34 507869
rect -96 506809 -62 507785
rect 62 506809 96 507785
rect -34 506725 34 506759
rect -34 506617 34 506651
rect -96 505591 -62 506567
rect 62 505591 96 506567
rect -34 505507 34 505541
rect -34 505399 34 505433
rect -96 504373 -62 505349
rect 62 504373 96 505349
rect -34 504289 34 504323
rect -34 504181 34 504215
rect -96 503155 -62 504131
rect 62 503155 96 504131
rect -34 503071 34 503105
rect -34 502963 34 502997
rect -96 501937 -62 502913
rect 62 501937 96 502913
rect -34 501853 34 501887
rect -34 501745 34 501779
rect -96 500719 -62 501695
rect 62 500719 96 501695
rect -34 500635 34 500669
rect -34 500527 34 500561
rect -96 499501 -62 500477
rect 62 499501 96 500477
rect -34 499417 34 499451
rect -34 499309 34 499343
rect -96 498283 -62 499259
rect 62 498283 96 499259
rect -34 498199 34 498233
rect -34 498091 34 498125
rect -96 497065 -62 498041
rect 62 497065 96 498041
rect -34 496981 34 497015
rect -34 496873 34 496907
rect -96 495847 -62 496823
rect 62 495847 96 496823
rect -34 495763 34 495797
rect -34 495655 34 495689
rect -96 494629 -62 495605
rect 62 494629 96 495605
rect -34 494545 34 494579
rect -34 494437 34 494471
rect -96 493411 -62 494387
rect 62 493411 96 494387
rect -34 493327 34 493361
rect -34 493219 34 493253
rect -96 492193 -62 493169
rect 62 492193 96 493169
rect -34 492109 34 492143
rect -34 492001 34 492035
rect -96 490975 -62 491951
rect 62 490975 96 491951
rect -34 490891 34 490925
rect -34 490783 34 490817
rect -96 489757 -62 490733
rect 62 489757 96 490733
rect -34 489673 34 489707
rect -34 489565 34 489599
rect -96 488539 -62 489515
rect 62 488539 96 489515
rect -34 488455 34 488489
rect -34 488347 34 488381
rect -96 487321 -62 488297
rect 62 487321 96 488297
rect -34 487237 34 487271
rect -34 487129 34 487163
rect -96 486103 -62 487079
rect 62 486103 96 487079
rect -34 486019 34 486053
rect -34 485911 34 485945
rect -96 484885 -62 485861
rect 62 484885 96 485861
rect -34 484801 34 484835
rect -34 484693 34 484727
rect -96 483667 -62 484643
rect 62 483667 96 484643
rect -34 483583 34 483617
rect -34 483475 34 483509
rect -96 482449 -62 483425
rect 62 482449 96 483425
rect -34 482365 34 482399
rect -34 482257 34 482291
rect -96 481231 -62 482207
rect 62 481231 96 482207
rect -34 481147 34 481181
rect -34 481039 34 481073
rect -96 480013 -62 480989
rect 62 480013 96 480989
rect -34 479929 34 479963
rect -34 479821 34 479855
rect -96 478795 -62 479771
rect 62 478795 96 479771
rect -34 478711 34 478745
rect -34 478603 34 478637
rect -96 477577 -62 478553
rect 62 477577 96 478553
rect -34 477493 34 477527
rect -34 477385 34 477419
rect -96 476359 -62 477335
rect 62 476359 96 477335
rect -34 476275 34 476309
rect -34 476167 34 476201
rect -96 475141 -62 476117
rect 62 475141 96 476117
rect -34 475057 34 475091
rect -34 474949 34 474983
rect -96 473923 -62 474899
rect 62 473923 96 474899
rect -34 473839 34 473873
rect -34 473731 34 473765
rect -96 472705 -62 473681
rect 62 472705 96 473681
rect -34 472621 34 472655
rect -34 472513 34 472547
rect -96 471487 -62 472463
rect 62 471487 96 472463
rect -34 471403 34 471437
rect -34 471295 34 471329
rect -96 470269 -62 471245
rect 62 470269 96 471245
rect -34 470185 34 470219
rect -34 470077 34 470111
rect -96 469051 -62 470027
rect 62 469051 96 470027
rect -34 468967 34 469001
rect -34 468859 34 468893
rect -96 467833 -62 468809
rect 62 467833 96 468809
rect -34 467749 34 467783
rect -34 467641 34 467675
rect -96 466615 -62 467591
rect 62 466615 96 467591
rect -34 466531 34 466565
rect -34 466423 34 466457
rect -96 465397 -62 466373
rect 62 465397 96 466373
rect -34 465313 34 465347
rect -34 465205 34 465239
rect -96 464179 -62 465155
rect 62 464179 96 465155
rect -34 464095 34 464129
rect -34 463987 34 464021
rect -96 462961 -62 463937
rect 62 462961 96 463937
rect -34 462877 34 462911
rect -34 462769 34 462803
rect -96 461743 -62 462719
rect 62 461743 96 462719
rect -34 461659 34 461693
rect -34 461551 34 461585
rect -96 460525 -62 461501
rect 62 460525 96 461501
rect -34 460441 34 460475
rect -34 460333 34 460367
rect -96 459307 -62 460283
rect 62 459307 96 460283
rect -34 459223 34 459257
rect -34 459115 34 459149
rect -96 458089 -62 459065
rect 62 458089 96 459065
rect -34 458005 34 458039
rect -34 457897 34 457931
rect -96 456871 -62 457847
rect 62 456871 96 457847
rect -34 456787 34 456821
rect -34 456679 34 456713
rect -96 455653 -62 456629
rect 62 455653 96 456629
rect -34 455569 34 455603
rect -34 455461 34 455495
rect -96 454435 -62 455411
rect 62 454435 96 455411
rect -34 454351 34 454385
rect -34 454243 34 454277
rect -96 453217 -62 454193
rect 62 453217 96 454193
rect -34 453133 34 453167
rect -34 453025 34 453059
rect -96 451999 -62 452975
rect 62 451999 96 452975
rect -34 451915 34 451949
rect -34 451807 34 451841
rect -96 450781 -62 451757
rect 62 450781 96 451757
rect -34 450697 34 450731
rect -34 450589 34 450623
rect -96 449563 -62 450539
rect 62 449563 96 450539
rect -34 449479 34 449513
rect -34 449371 34 449405
rect -96 448345 -62 449321
rect 62 448345 96 449321
rect -34 448261 34 448295
rect -34 448153 34 448187
rect -96 447127 -62 448103
rect 62 447127 96 448103
rect -34 447043 34 447077
rect -34 446935 34 446969
rect -96 445909 -62 446885
rect 62 445909 96 446885
rect -34 445825 34 445859
rect -34 445717 34 445751
rect -96 444691 -62 445667
rect 62 444691 96 445667
rect -34 444607 34 444641
rect -34 444499 34 444533
rect -96 443473 -62 444449
rect 62 443473 96 444449
rect -34 443389 34 443423
rect -34 443281 34 443315
rect -96 442255 -62 443231
rect 62 442255 96 443231
rect -34 442171 34 442205
rect -34 442063 34 442097
rect -96 441037 -62 442013
rect 62 441037 96 442013
rect -34 440953 34 440987
rect -34 440845 34 440879
rect -96 439819 -62 440795
rect 62 439819 96 440795
rect -34 439735 34 439769
rect -34 439627 34 439661
rect -96 438601 -62 439577
rect 62 438601 96 439577
rect -34 438517 34 438551
rect -34 438409 34 438443
rect -96 437383 -62 438359
rect 62 437383 96 438359
rect -34 437299 34 437333
rect -34 437191 34 437225
rect -96 436165 -62 437141
rect 62 436165 96 437141
rect -34 436081 34 436115
rect -34 435973 34 436007
rect -96 434947 -62 435923
rect 62 434947 96 435923
rect -34 434863 34 434897
rect -34 434755 34 434789
rect -96 433729 -62 434705
rect 62 433729 96 434705
rect -34 433645 34 433679
rect -34 433537 34 433571
rect -96 432511 -62 433487
rect 62 432511 96 433487
rect -34 432427 34 432461
rect -34 432319 34 432353
rect -96 431293 -62 432269
rect 62 431293 96 432269
rect -34 431209 34 431243
rect -34 431101 34 431135
rect -96 430075 -62 431051
rect 62 430075 96 431051
rect -34 429991 34 430025
rect -34 429883 34 429917
rect -96 428857 -62 429833
rect 62 428857 96 429833
rect -34 428773 34 428807
rect -34 428665 34 428699
rect -96 427639 -62 428615
rect 62 427639 96 428615
rect -34 427555 34 427589
rect -34 427447 34 427481
rect -96 426421 -62 427397
rect 62 426421 96 427397
rect -34 426337 34 426371
rect -34 426229 34 426263
rect -96 425203 -62 426179
rect 62 425203 96 426179
rect -34 425119 34 425153
rect -34 425011 34 425045
rect -96 423985 -62 424961
rect 62 423985 96 424961
rect -34 423901 34 423935
rect -34 423793 34 423827
rect -96 422767 -62 423743
rect 62 422767 96 423743
rect -34 422683 34 422717
rect -34 422575 34 422609
rect -96 421549 -62 422525
rect 62 421549 96 422525
rect -34 421465 34 421499
rect -34 421357 34 421391
rect -96 420331 -62 421307
rect 62 420331 96 421307
rect -34 420247 34 420281
rect -34 420139 34 420173
rect -96 419113 -62 420089
rect 62 419113 96 420089
rect -34 419029 34 419063
rect -34 418921 34 418955
rect -96 417895 -62 418871
rect 62 417895 96 418871
rect -34 417811 34 417845
rect -34 417703 34 417737
rect -96 416677 -62 417653
rect 62 416677 96 417653
rect -34 416593 34 416627
rect -34 416485 34 416519
rect -96 415459 -62 416435
rect 62 415459 96 416435
rect -34 415375 34 415409
rect -34 415267 34 415301
rect -96 414241 -62 415217
rect 62 414241 96 415217
rect -34 414157 34 414191
rect -34 414049 34 414083
rect -96 413023 -62 413999
rect 62 413023 96 413999
rect -34 412939 34 412973
rect -34 412831 34 412865
rect -96 411805 -62 412781
rect 62 411805 96 412781
rect -34 411721 34 411755
rect -34 411613 34 411647
rect -96 410587 -62 411563
rect 62 410587 96 411563
rect -34 410503 34 410537
rect -34 410395 34 410429
rect -96 409369 -62 410345
rect 62 409369 96 410345
rect -34 409285 34 409319
rect -34 409177 34 409211
rect -96 408151 -62 409127
rect 62 408151 96 409127
rect -34 408067 34 408101
rect -34 407959 34 407993
rect -96 406933 -62 407909
rect 62 406933 96 407909
rect -34 406849 34 406883
rect -34 406741 34 406775
rect -96 405715 -62 406691
rect 62 405715 96 406691
rect -34 405631 34 405665
rect -34 405523 34 405557
rect -96 404497 -62 405473
rect 62 404497 96 405473
rect -34 404413 34 404447
rect -34 404305 34 404339
rect -96 403279 -62 404255
rect 62 403279 96 404255
rect -34 403195 34 403229
rect -34 403087 34 403121
rect -96 402061 -62 403037
rect 62 402061 96 403037
rect -34 401977 34 402011
rect -34 401869 34 401903
rect -96 400843 -62 401819
rect 62 400843 96 401819
rect -34 400759 34 400793
rect -34 400651 34 400685
rect -96 399625 -62 400601
rect 62 399625 96 400601
rect -34 399541 34 399575
rect -34 399433 34 399467
rect -96 398407 -62 399383
rect 62 398407 96 399383
rect -34 398323 34 398357
rect -34 398215 34 398249
rect -96 397189 -62 398165
rect 62 397189 96 398165
rect -34 397105 34 397139
rect -34 396997 34 397031
rect -96 395971 -62 396947
rect 62 395971 96 396947
rect -34 395887 34 395921
rect -34 395779 34 395813
rect -96 394753 -62 395729
rect 62 394753 96 395729
rect -34 394669 34 394703
rect -34 394561 34 394595
rect -96 393535 -62 394511
rect 62 393535 96 394511
rect -34 393451 34 393485
rect -34 393343 34 393377
rect -96 392317 -62 393293
rect 62 392317 96 393293
rect -34 392233 34 392267
rect -34 392125 34 392159
rect -96 391099 -62 392075
rect 62 391099 96 392075
rect -34 391015 34 391049
rect -34 390907 34 390941
rect -96 389881 -62 390857
rect 62 389881 96 390857
rect -34 389797 34 389831
rect -34 389689 34 389723
rect -96 388663 -62 389639
rect 62 388663 96 389639
rect -34 388579 34 388613
rect -34 388471 34 388505
rect -96 387445 -62 388421
rect 62 387445 96 388421
rect -34 387361 34 387395
rect -34 387253 34 387287
rect -96 386227 -62 387203
rect 62 386227 96 387203
rect -34 386143 34 386177
rect -34 386035 34 386069
rect -96 385009 -62 385985
rect 62 385009 96 385985
rect -34 384925 34 384959
rect -34 384817 34 384851
rect -96 383791 -62 384767
rect 62 383791 96 384767
rect -34 383707 34 383741
rect -34 383599 34 383633
rect -96 382573 -62 383549
rect 62 382573 96 383549
rect -34 382489 34 382523
rect -34 382381 34 382415
rect -96 381355 -62 382331
rect 62 381355 96 382331
rect -34 381271 34 381305
rect -34 381163 34 381197
rect -96 380137 -62 381113
rect 62 380137 96 381113
rect -34 380053 34 380087
rect -34 379945 34 379979
rect -96 378919 -62 379895
rect 62 378919 96 379895
rect -34 378835 34 378869
rect -34 378727 34 378761
rect -96 377701 -62 378677
rect 62 377701 96 378677
rect -34 377617 34 377651
rect -34 377509 34 377543
rect -96 376483 -62 377459
rect 62 376483 96 377459
rect -34 376399 34 376433
rect -34 376291 34 376325
rect -96 375265 -62 376241
rect 62 375265 96 376241
rect -34 375181 34 375215
rect -34 375073 34 375107
rect -96 374047 -62 375023
rect 62 374047 96 375023
rect -34 373963 34 373997
rect -34 373855 34 373889
rect -96 372829 -62 373805
rect 62 372829 96 373805
rect -34 372745 34 372779
rect -34 372637 34 372671
rect -96 371611 -62 372587
rect 62 371611 96 372587
rect -34 371527 34 371561
rect -34 371419 34 371453
rect -96 370393 -62 371369
rect 62 370393 96 371369
rect -34 370309 34 370343
rect -34 370201 34 370235
rect -96 369175 -62 370151
rect 62 369175 96 370151
rect -34 369091 34 369125
rect -34 368983 34 369017
rect -96 367957 -62 368933
rect 62 367957 96 368933
rect -34 367873 34 367907
rect -34 367765 34 367799
rect -96 366739 -62 367715
rect 62 366739 96 367715
rect -34 366655 34 366689
rect -34 366547 34 366581
rect -96 365521 -62 366497
rect 62 365521 96 366497
rect -34 365437 34 365471
rect -34 365329 34 365363
rect -96 364303 -62 365279
rect 62 364303 96 365279
rect -34 364219 34 364253
rect -34 364111 34 364145
rect -96 363085 -62 364061
rect 62 363085 96 364061
rect -34 363001 34 363035
rect -34 362893 34 362927
rect -96 361867 -62 362843
rect 62 361867 96 362843
rect -34 361783 34 361817
rect -34 361675 34 361709
rect -96 360649 -62 361625
rect 62 360649 96 361625
rect -34 360565 34 360599
rect -34 360457 34 360491
rect -96 359431 -62 360407
rect 62 359431 96 360407
rect -34 359347 34 359381
rect -34 359239 34 359273
rect -96 358213 -62 359189
rect 62 358213 96 359189
rect -34 358129 34 358163
rect -34 358021 34 358055
rect -96 356995 -62 357971
rect 62 356995 96 357971
rect -34 356911 34 356945
rect -34 356803 34 356837
rect -96 355777 -62 356753
rect 62 355777 96 356753
rect -34 355693 34 355727
rect -34 355585 34 355619
rect -96 354559 -62 355535
rect 62 354559 96 355535
rect -34 354475 34 354509
rect -34 354367 34 354401
rect -96 353341 -62 354317
rect 62 353341 96 354317
rect -34 353257 34 353291
rect -34 353149 34 353183
rect -96 352123 -62 353099
rect 62 352123 96 353099
rect -34 352039 34 352073
rect -34 351931 34 351965
rect -96 350905 -62 351881
rect 62 350905 96 351881
rect -34 350821 34 350855
rect -34 350713 34 350747
rect -96 349687 -62 350663
rect 62 349687 96 350663
rect -34 349603 34 349637
rect -34 349495 34 349529
rect -96 348469 -62 349445
rect 62 348469 96 349445
rect -34 348385 34 348419
rect -34 348277 34 348311
rect -96 347251 -62 348227
rect 62 347251 96 348227
rect -34 347167 34 347201
rect -34 347059 34 347093
rect -96 346033 -62 347009
rect 62 346033 96 347009
rect -34 345949 34 345983
rect -34 345841 34 345875
rect -96 344815 -62 345791
rect 62 344815 96 345791
rect -34 344731 34 344765
rect -34 344623 34 344657
rect -96 343597 -62 344573
rect 62 343597 96 344573
rect -34 343513 34 343547
rect -34 343405 34 343439
rect -96 342379 -62 343355
rect 62 342379 96 343355
rect -34 342295 34 342329
rect -34 342187 34 342221
rect -96 341161 -62 342137
rect 62 341161 96 342137
rect -34 341077 34 341111
rect -34 340969 34 341003
rect -96 339943 -62 340919
rect 62 339943 96 340919
rect -34 339859 34 339893
rect -34 339751 34 339785
rect -96 338725 -62 339701
rect 62 338725 96 339701
rect -34 338641 34 338675
rect -34 338533 34 338567
rect -96 337507 -62 338483
rect 62 337507 96 338483
rect -34 337423 34 337457
rect -34 337315 34 337349
rect -96 336289 -62 337265
rect 62 336289 96 337265
rect -34 336205 34 336239
rect -34 336097 34 336131
rect -96 335071 -62 336047
rect 62 335071 96 336047
rect -34 334987 34 335021
rect -34 334879 34 334913
rect -96 333853 -62 334829
rect 62 333853 96 334829
rect -34 333769 34 333803
rect -34 333661 34 333695
rect -96 332635 -62 333611
rect 62 332635 96 333611
rect -34 332551 34 332585
rect -34 332443 34 332477
rect -96 331417 -62 332393
rect 62 331417 96 332393
rect -34 331333 34 331367
rect -34 331225 34 331259
rect -96 330199 -62 331175
rect 62 330199 96 331175
rect -34 330115 34 330149
rect -34 330007 34 330041
rect -96 328981 -62 329957
rect 62 328981 96 329957
rect -34 328897 34 328931
rect -34 328789 34 328823
rect -96 327763 -62 328739
rect 62 327763 96 328739
rect -34 327679 34 327713
rect -34 327571 34 327605
rect -96 326545 -62 327521
rect 62 326545 96 327521
rect -34 326461 34 326495
rect -34 326353 34 326387
rect -96 325327 -62 326303
rect 62 325327 96 326303
rect -34 325243 34 325277
rect -34 325135 34 325169
rect -96 324109 -62 325085
rect 62 324109 96 325085
rect -34 324025 34 324059
rect -34 323917 34 323951
rect -96 322891 -62 323867
rect 62 322891 96 323867
rect -34 322807 34 322841
rect -34 322699 34 322733
rect -96 321673 -62 322649
rect 62 321673 96 322649
rect -34 321589 34 321623
rect -34 321481 34 321515
rect -96 320455 -62 321431
rect 62 320455 96 321431
rect -34 320371 34 320405
rect -34 320263 34 320297
rect -96 319237 -62 320213
rect 62 319237 96 320213
rect -34 319153 34 319187
rect -34 319045 34 319079
rect -96 318019 -62 318995
rect 62 318019 96 318995
rect -34 317935 34 317969
rect -34 317827 34 317861
rect -96 316801 -62 317777
rect 62 316801 96 317777
rect -34 316717 34 316751
rect -34 316609 34 316643
rect -96 315583 -62 316559
rect 62 315583 96 316559
rect -34 315499 34 315533
rect -34 315391 34 315425
rect -96 314365 -62 315341
rect 62 314365 96 315341
rect -34 314281 34 314315
rect -34 314173 34 314207
rect -96 313147 -62 314123
rect 62 313147 96 314123
rect -34 313063 34 313097
rect -34 312955 34 312989
rect -96 311929 -62 312905
rect 62 311929 96 312905
rect -34 311845 34 311879
rect -34 311737 34 311771
rect -96 310711 -62 311687
rect 62 310711 96 311687
rect -34 310627 34 310661
rect -34 310519 34 310553
rect -96 309493 -62 310469
rect 62 309493 96 310469
rect -34 309409 34 309443
rect -34 309301 34 309335
rect -96 308275 -62 309251
rect 62 308275 96 309251
rect -34 308191 34 308225
rect -34 308083 34 308117
rect -96 307057 -62 308033
rect 62 307057 96 308033
rect -34 306973 34 307007
rect -34 306865 34 306899
rect -96 305839 -62 306815
rect 62 305839 96 306815
rect -34 305755 34 305789
rect -34 305647 34 305681
rect -96 304621 -62 305597
rect 62 304621 96 305597
rect -34 304537 34 304571
rect -34 304429 34 304463
rect -96 303403 -62 304379
rect 62 303403 96 304379
rect -34 303319 34 303353
rect -34 303211 34 303245
rect -96 302185 -62 303161
rect 62 302185 96 303161
rect -34 302101 34 302135
rect -34 301993 34 302027
rect -96 300967 -62 301943
rect 62 300967 96 301943
rect -34 300883 34 300917
rect -34 300775 34 300809
rect -96 299749 -62 300725
rect 62 299749 96 300725
rect -34 299665 34 299699
rect -34 299557 34 299591
rect -96 298531 -62 299507
rect 62 298531 96 299507
rect -34 298447 34 298481
rect -34 298339 34 298373
rect -96 297313 -62 298289
rect 62 297313 96 298289
rect -34 297229 34 297263
rect -34 297121 34 297155
rect -96 296095 -62 297071
rect 62 296095 96 297071
rect -34 296011 34 296045
rect -34 295903 34 295937
rect -96 294877 -62 295853
rect 62 294877 96 295853
rect -34 294793 34 294827
rect -34 294685 34 294719
rect -96 293659 -62 294635
rect 62 293659 96 294635
rect -34 293575 34 293609
rect -34 293467 34 293501
rect -96 292441 -62 293417
rect 62 292441 96 293417
rect -34 292357 34 292391
rect -34 292249 34 292283
rect -96 291223 -62 292199
rect 62 291223 96 292199
rect -34 291139 34 291173
rect -34 291031 34 291065
rect -96 290005 -62 290981
rect 62 290005 96 290981
rect -34 289921 34 289955
rect -34 289813 34 289847
rect -96 288787 -62 289763
rect 62 288787 96 289763
rect -34 288703 34 288737
rect -34 288595 34 288629
rect -96 287569 -62 288545
rect 62 287569 96 288545
rect -34 287485 34 287519
rect -34 287377 34 287411
rect -96 286351 -62 287327
rect 62 286351 96 287327
rect -34 286267 34 286301
rect -34 286159 34 286193
rect -96 285133 -62 286109
rect 62 285133 96 286109
rect -34 285049 34 285083
rect -34 284941 34 284975
rect -96 283915 -62 284891
rect 62 283915 96 284891
rect -34 283831 34 283865
rect -34 283723 34 283757
rect -96 282697 -62 283673
rect 62 282697 96 283673
rect -34 282613 34 282647
rect -34 282505 34 282539
rect -96 281479 -62 282455
rect 62 281479 96 282455
rect -34 281395 34 281429
rect -34 281287 34 281321
rect -96 280261 -62 281237
rect 62 280261 96 281237
rect -34 280177 34 280211
rect -34 280069 34 280103
rect -96 279043 -62 280019
rect 62 279043 96 280019
rect -34 278959 34 278993
rect -34 278851 34 278885
rect -96 277825 -62 278801
rect 62 277825 96 278801
rect -34 277741 34 277775
rect -34 277633 34 277667
rect -96 276607 -62 277583
rect 62 276607 96 277583
rect -34 276523 34 276557
rect -34 276415 34 276449
rect -96 275389 -62 276365
rect 62 275389 96 276365
rect -34 275305 34 275339
rect -34 275197 34 275231
rect -96 274171 -62 275147
rect 62 274171 96 275147
rect -34 274087 34 274121
rect -34 273979 34 274013
rect -96 272953 -62 273929
rect 62 272953 96 273929
rect -34 272869 34 272903
rect -34 272761 34 272795
rect -96 271735 -62 272711
rect 62 271735 96 272711
rect -34 271651 34 271685
rect -34 271543 34 271577
rect -96 270517 -62 271493
rect 62 270517 96 271493
rect -34 270433 34 270467
rect -34 270325 34 270359
rect -96 269299 -62 270275
rect 62 269299 96 270275
rect -34 269215 34 269249
rect -34 269107 34 269141
rect -96 268081 -62 269057
rect 62 268081 96 269057
rect -34 267997 34 268031
rect -34 267889 34 267923
rect -96 266863 -62 267839
rect 62 266863 96 267839
rect -34 266779 34 266813
rect -34 266671 34 266705
rect -96 265645 -62 266621
rect 62 265645 96 266621
rect -34 265561 34 265595
rect -34 265453 34 265487
rect -96 264427 -62 265403
rect 62 264427 96 265403
rect -34 264343 34 264377
rect -34 264235 34 264269
rect -96 263209 -62 264185
rect 62 263209 96 264185
rect -34 263125 34 263159
rect -34 263017 34 263051
rect -96 261991 -62 262967
rect 62 261991 96 262967
rect -34 261907 34 261941
rect -34 261799 34 261833
rect -96 260773 -62 261749
rect 62 260773 96 261749
rect -34 260689 34 260723
rect -34 260581 34 260615
rect -96 259555 -62 260531
rect 62 259555 96 260531
rect -34 259471 34 259505
rect -34 259363 34 259397
rect -96 258337 -62 259313
rect 62 258337 96 259313
rect -34 258253 34 258287
rect -34 258145 34 258179
rect -96 257119 -62 258095
rect 62 257119 96 258095
rect -34 257035 34 257069
rect -34 256927 34 256961
rect -96 255901 -62 256877
rect 62 255901 96 256877
rect -34 255817 34 255851
rect -34 255709 34 255743
rect -96 254683 -62 255659
rect 62 254683 96 255659
rect -34 254599 34 254633
rect -34 254491 34 254525
rect -96 253465 -62 254441
rect 62 253465 96 254441
rect -34 253381 34 253415
rect -34 253273 34 253307
rect -96 252247 -62 253223
rect 62 252247 96 253223
rect -34 252163 34 252197
rect -34 252055 34 252089
rect -96 251029 -62 252005
rect 62 251029 96 252005
rect -34 250945 34 250979
rect -34 250837 34 250871
rect -96 249811 -62 250787
rect 62 249811 96 250787
rect -34 249727 34 249761
rect -34 249619 34 249653
rect -96 248593 -62 249569
rect 62 248593 96 249569
rect -34 248509 34 248543
rect -34 248401 34 248435
rect -96 247375 -62 248351
rect 62 247375 96 248351
rect -34 247291 34 247325
rect -34 247183 34 247217
rect -96 246157 -62 247133
rect 62 246157 96 247133
rect -34 246073 34 246107
rect -34 245965 34 245999
rect -96 244939 -62 245915
rect 62 244939 96 245915
rect -34 244855 34 244889
rect -34 244747 34 244781
rect -96 243721 -62 244697
rect 62 243721 96 244697
rect -34 243637 34 243671
rect -34 243529 34 243563
rect -96 242503 -62 243479
rect 62 242503 96 243479
rect -34 242419 34 242453
rect -34 242311 34 242345
rect -96 241285 -62 242261
rect 62 241285 96 242261
rect -34 241201 34 241235
rect -34 241093 34 241127
rect -96 240067 -62 241043
rect 62 240067 96 241043
rect -34 239983 34 240017
rect -34 239875 34 239909
rect -96 238849 -62 239825
rect 62 238849 96 239825
rect -34 238765 34 238799
rect -34 238657 34 238691
rect -96 237631 -62 238607
rect 62 237631 96 238607
rect -34 237547 34 237581
rect -34 237439 34 237473
rect -96 236413 -62 237389
rect 62 236413 96 237389
rect -34 236329 34 236363
rect -34 236221 34 236255
rect -96 235195 -62 236171
rect 62 235195 96 236171
rect -34 235111 34 235145
rect -34 235003 34 235037
rect -96 233977 -62 234953
rect 62 233977 96 234953
rect -34 233893 34 233927
rect -34 233785 34 233819
rect -96 232759 -62 233735
rect 62 232759 96 233735
rect -34 232675 34 232709
rect -34 232567 34 232601
rect -96 231541 -62 232517
rect 62 231541 96 232517
rect -34 231457 34 231491
rect -34 231349 34 231383
rect -96 230323 -62 231299
rect 62 230323 96 231299
rect -34 230239 34 230273
rect -34 230131 34 230165
rect -96 229105 -62 230081
rect 62 229105 96 230081
rect -34 229021 34 229055
rect -34 228913 34 228947
rect -96 227887 -62 228863
rect 62 227887 96 228863
rect -34 227803 34 227837
rect -34 227695 34 227729
rect -96 226669 -62 227645
rect 62 226669 96 227645
rect -34 226585 34 226619
rect -34 226477 34 226511
rect -96 225451 -62 226427
rect 62 225451 96 226427
rect -34 225367 34 225401
rect -34 225259 34 225293
rect -96 224233 -62 225209
rect 62 224233 96 225209
rect -34 224149 34 224183
rect -34 224041 34 224075
rect -96 223015 -62 223991
rect 62 223015 96 223991
rect -34 222931 34 222965
rect -34 222823 34 222857
rect -96 221797 -62 222773
rect 62 221797 96 222773
rect -34 221713 34 221747
rect -34 221605 34 221639
rect -96 220579 -62 221555
rect 62 220579 96 221555
rect -34 220495 34 220529
rect -34 220387 34 220421
rect -96 219361 -62 220337
rect 62 219361 96 220337
rect -34 219277 34 219311
rect -34 219169 34 219203
rect -96 218143 -62 219119
rect 62 218143 96 219119
rect -34 218059 34 218093
rect -34 217951 34 217985
rect -96 216925 -62 217901
rect 62 216925 96 217901
rect -34 216841 34 216875
rect -34 216733 34 216767
rect -96 215707 -62 216683
rect 62 215707 96 216683
rect -34 215623 34 215657
rect -34 215515 34 215549
rect -96 214489 -62 215465
rect 62 214489 96 215465
rect -34 214405 34 214439
rect -34 214297 34 214331
rect -96 213271 -62 214247
rect 62 213271 96 214247
rect -34 213187 34 213221
rect -34 213079 34 213113
rect -96 212053 -62 213029
rect 62 212053 96 213029
rect -34 211969 34 212003
rect -34 211861 34 211895
rect -96 210835 -62 211811
rect 62 210835 96 211811
rect -34 210751 34 210785
rect -34 210643 34 210677
rect -96 209617 -62 210593
rect 62 209617 96 210593
rect -34 209533 34 209567
rect -34 209425 34 209459
rect -96 208399 -62 209375
rect 62 208399 96 209375
rect -34 208315 34 208349
rect -34 208207 34 208241
rect -96 207181 -62 208157
rect 62 207181 96 208157
rect -34 207097 34 207131
rect -34 206989 34 207023
rect -96 205963 -62 206939
rect 62 205963 96 206939
rect -34 205879 34 205913
rect -34 205771 34 205805
rect -96 204745 -62 205721
rect 62 204745 96 205721
rect -34 204661 34 204695
rect -34 204553 34 204587
rect -96 203527 -62 204503
rect 62 203527 96 204503
rect -34 203443 34 203477
rect -34 203335 34 203369
rect -96 202309 -62 203285
rect 62 202309 96 203285
rect -34 202225 34 202259
rect -34 202117 34 202151
rect -96 201091 -62 202067
rect 62 201091 96 202067
rect -34 201007 34 201041
rect -34 200899 34 200933
rect -96 199873 -62 200849
rect 62 199873 96 200849
rect -34 199789 34 199823
rect -34 199681 34 199715
rect -96 198655 -62 199631
rect 62 198655 96 199631
rect -34 198571 34 198605
rect -34 198463 34 198497
rect -96 197437 -62 198413
rect 62 197437 96 198413
rect -34 197353 34 197387
rect -34 197245 34 197279
rect -96 196219 -62 197195
rect 62 196219 96 197195
rect -34 196135 34 196169
rect -34 196027 34 196061
rect -96 195001 -62 195977
rect 62 195001 96 195977
rect -34 194917 34 194951
rect -34 194809 34 194843
rect -96 193783 -62 194759
rect 62 193783 96 194759
rect -34 193699 34 193733
rect -34 193591 34 193625
rect -96 192565 -62 193541
rect 62 192565 96 193541
rect -34 192481 34 192515
rect -34 192373 34 192407
rect -96 191347 -62 192323
rect 62 191347 96 192323
rect -34 191263 34 191297
rect -34 191155 34 191189
rect -96 190129 -62 191105
rect 62 190129 96 191105
rect -34 190045 34 190079
rect -34 189937 34 189971
rect -96 188911 -62 189887
rect 62 188911 96 189887
rect -34 188827 34 188861
rect -34 188719 34 188753
rect -96 187693 -62 188669
rect 62 187693 96 188669
rect -34 187609 34 187643
rect -34 187501 34 187535
rect -96 186475 -62 187451
rect 62 186475 96 187451
rect -34 186391 34 186425
rect -34 186283 34 186317
rect -96 185257 -62 186233
rect 62 185257 96 186233
rect -34 185173 34 185207
rect -34 185065 34 185099
rect -96 184039 -62 185015
rect 62 184039 96 185015
rect -34 183955 34 183989
rect -34 183847 34 183881
rect -96 182821 -62 183797
rect 62 182821 96 183797
rect -34 182737 34 182771
rect -34 182629 34 182663
rect -96 181603 -62 182579
rect 62 181603 96 182579
rect -34 181519 34 181553
rect -34 181411 34 181445
rect -96 180385 -62 181361
rect 62 180385 96 181361
rect -34 180301 34 180335
rect -34 180193 34 180227
rect -96 179167 -62 180143
rect 62 179167 96 180143
rect -34 179083 34 179117
rect -34 178975 34 179009
rect -96 177949 -62 178925
rect 62 177949 96 178925
rect -34 177865 34 177899
rect -34 177757 34 177791
rect -96 176731 -62 177707
rect 62 176731 96 177707
rect -34 176647 34 176681
rect -34 176539 34 176573
rect -96 175513 -62 176489
rect 62 175513 96 176489
rect -34 175429 34 175463
rect -34 175321 34 175355
rect -96 174295 -62 175271
rect 62 174295 96 175271
rect -34 174211 34 174245
rect -34 174103 34 174137
rect -96 173077 -62 174053
rect 62 173077 96 174053
rect -34 172993 34 173027
rect -34 172885 34 172919
rect -96 171859 -62 172835
rect 62 171859 96 172835
rect -34 171775 34 171809
rect -34 171667 34 171701
rect -96 170641 -62 171617
rect 62 170641 96 171617
rect -34 170557 34 170591
rect -34 170449 34 170483
rect -96 169423 -62 170399
rect 62 169423 96 170399
rect -34 169339 34 169373
rect -34 169231 34 169265
rect -96 168205 -62 169181
rect 62 168205 96 169181
rect -34 168121 34 168155
rect -34 168013 34 168047
rect -96 166987 -62 167963
rect 62 166987 96 167963
rect -34 166903 34 166937
rect -34 166795 34 166829
rect -96 165769 -62 166745
rect 62 165769 96 166745
rect -34 165685 34 165719
rect -34 165577 34 165611
rect -96 164551 -62 165527
rect 62 164551 96 165527
rect -34 164467 34 164501
rect -34 164359 34 164393
rect -96 163333 -62 164309
rect 62 163333 96 164309
rect -34 163249 34 163283
rect -34 163141 34 163175
rect -96 162115 -62 163091
rect 62 162115 96 163091
rect -34 162031 34 162065
rect -34 161923 34 161957
rect -96 160897 -62 161873
rect 62 160897 96 161873
rect -34 160813 34 160847
rect -34 160705 34 160739
rect -96 159679 -62 160655
rect 62 159679 96 160655
rect -34 159595 34 159629
rect -34 159487 34 159521
rect -96 158461 -62 159437
rect 62 158461 96 159437
rect -34 158377 34 158411
rect -34 158269 34 158303
rect -96 157243 -62 158219
rect 62 157243 96 158219
rect -34 157159 34 157193
rect -34 157051 34 157085
rect -96 156025 -62 157001
rect 62 156025 96 157001
rect -34 155941 34 155975
rect -34 155833 34 155867
rect -96 154807 -62 155783
rect 62 154807 96 155783
rect -34 154723 34 154757
rect -34 154615 34 154649
rect -96 153589 -62 154565
rect 62 153589 96 154565
rect -34 153505 34 153539
rect -34 153397 34 153431
rect -96 152371 -62 153347
rect 62 152371 96 153347
rect -34 152287 34 152321
rect -34 152179 34 152213
rect -96 151153 -62 152129
rect 62 151153 96 152129
rect -34 151069 34 151103
rect -34 150961 34 150995
rect -96 149935 -62 150911
rect 62 149935 96 150911
rect -34 149851 34 149885
rect -34 149743 34 149777
rect -96 148717 -62 149693
rect 62 148717 96 149693
rect -34 148633 34 148667
rect -34 148525 34 148559
rect -96 147499 -62 148475
rect 62 147499 96 148475
rect -34 147415 34 147449
rect -34 147307 34 147341
rect -96 146281 -62 147257
rect 62 146281 96 147257
rect -34 146197 34 146231
rect -34 146089 34 146123
rect -96 145063 -62 146039
rect 62 145063 96 146039
rect -34 144979 34 145013
rect -34 144871 34 144905
rect -96 143845 -62 144821
rect 62 143845 96 144821
rect -34 143761 34 143795
rect -34 143653 34 143687
rect -96 142627 -62 143603
rect 62 142627 96 143603
rect -34 142543 34 142577
rect -34 142435 34 142469
rect -96 141409 -62 142385
rect 62 141409 96 142385
rect -34 141325 34 141359
rect -34 141217 34 141251
rect -96 140191 -62 141167
rect 62 140191 96 141167
rect -34 140107 34 140141
rect -34 139999 34 140033
rect -96 138973 -62 139949
rect 62 138973 96 139949
rect -34 138889 34 138923
rect -34 138781 34 138815
rect -96 137755 -62 138731
rect 62 137755 96 138731
rect -34 137671 34 137705
rect -34 137563 34 137597
rect -96 136537 -62 137513
rect 62 136537 96 137513
rect -34 136453 34 136487
rect -34 136345 34 136379
rect -96 135319 -62 136295
rect 62 135319 96 136295
rect -34 135235 34 135269
rect -34 135127 34 135161
rect -96 134101 -62 135077
rect 62 134101 96 135077
rect -34 134017 34 134051
rect -34 133909 34 133943
rect -96 132883 -62 133859
rect 62 132883 96 133859
rect -34 132799 34 132833
rect -34 132691 34 132725
rect -96 131665 -62 132641
rect 62 131665 96 132641
rect -34 131581 34 131615
rect -34 131473 34 131507
rect -96 130447 -62 131423
rect 62 130447 96 131423
rect -34 130363 34 130397
rect -34 130255 34 130289
rect -96 129229 -62 130205
rect 62 129229 96 130205
rect -34 129145 34 129179
rect -34 129037 34 129071
rect -96 128011 -62 128987
rect 62 128011 96 128987
rect -34 127927 34 127961
rect -34 127819 34 127853
rect -96 126793 -62 127769
rect 62 126793 96 127769
rect -34 126709 34 126743
rect -34 126601 34 126635
rect -96 125575 -62 126551
rect 62 125575 96 126551
rect -34 125491 34 125525
rect -34 125383 34 125417
rect -96 124357 -62 125333
rect 62 124357 96 125333
rect -34 124273 34 124307
rect -34 124165 34 124199
rect -96 123139 -62 124115
rect 62 123139 96 124115
rect -34 123055 34 123089
rect -34 122947 34 122981
rect -96 121921 -62 122897
rect 62 121921 96 122897
rect -34 121837 34 121871
rect -34 121729 34 121763
rect -96 120703 -62 121679
rect 62 120703 96 121679
rect -34 120619 34 120653
rect -34 120511 34 120545
rect -96 119485 -62 120461
rect 62 119485 96 120461
rect -34 119401 34 119435
rect -34 119293 34 119327
rect -96 118267 -62 119243
rect 62 118267 96 119243
rect -34 118183 34 118217
rect -34 118075 34 118109
rect -96 117049 -62 118025
rect 62 117049 96 118025
rect -34 116965 34 116999
rect -34 116857 34 116891
rect -96 115831 -62 116807
rect 62 115831 96 116807
rect -34 115747 34 115781
rect -34 115639 34 115673
rect -96 114613 -62 115589
rect 62 114613 96 115589
rect -34 114529 34 114563
rect -34 114421 34 114455
rect -96 113395 -62 114371
rect 62 113395 96 114371
rect -34 113311 34 113345
rect -34 113203 34 113237
rect -96 112177 -62 113153
rect 62 112177 96 113153
rect -34 112093 34 112127
rect -34 111985 34 112019
rect -96 110959 -62 111935
rect 62 110959 96 111935
rect -34 110875 34 110909
rect -34 110767 34 110801
rect -96 109741 -62 110717
rect 62 109741 96 110717
rect -34 109657 34 109691
rect -34 109549 34 109583
rect -96 108523 -62 109499
rect 62 108523 96 109499
rect -34 108439 34 108473
rect -34 108331 34 108365
rect -96 107305 -62 108281
rect 62 107305 96 108281
rect -34 107221 34 107255
rect -34 107113 34 107147
rect -96 106087 -62 107063
rect 62 106087 96 107063
rect -34 106003 34 106037
rect -34 105895 34 105929
rect -96 104869 -62 105845
rect 62 104869 96 105845
rect -34 104785 34 104819
rect -34 104677 34 104711
rect -96 103651 -62 104627
rect 62 103651 96 104627
rect -34 103567 34 103601
rect -34 103459 34 103493
rect -96 102433 -62 103409
rect 62 102433 96 103409
rect -34 102349 34 102383
rect -34 102241 34 102275
rect -96 101215 -62 102191
rect 62 101215 96 102191
rect -34 101131 34 101165
rect -34 101023 34 101057
rect -96 99997 -62 100973
rect 62 99997 96 100973
rect -34 99913 34 99947
rect -34 99805 34 99839
rect -96 98779 -62 99755
rect 62 98779 96 99755
rect -34 98695 34 98729
rect -34 98587 34 98621
rect -96 97561 -62 98537
rect 62 97561 96 98537
rect -34 97477 34 97511
rect -34 97369 34 97403
rect -96 96343 -62 97319
rect 62 96343 96 97319
rect -34 96259 34 96293
rect -34 96151 34 96185
rect -96 95125 -62 96101
rect 62 95125 96 96101
rect -34 95041 34 95075
rect -34 94933 34 94967
rect -96 93907 -62 94883
rect 62 93907 96 94883
rect -34 93823 34 93857
rect -34 93715 34 93749
rect -96 92689 -62 93665
rect 62 92689 96 93665
rect -34 92605 34 92639
rect -34 92497 34 92531
rect -96 91471 -62 92447
rect 62 91471 96 92447
rect -34 91387 34 91421
rect -34 91279 34 91313
rect -96 90253 -62 91229
rect 62 90253 96 91229
rect -34 90169 34 90203
rect -34 90061 34 90095
rect -96 89035 -62 90011
rect 62 89035 96 90011
rect -34 88951 34 88985
rect -34 88843 34 88877
rect -96 87817 -62 88793
rect 62 87817 96 88793
rect -34 87733 34 87767
rect -34 87625 34 87659
rect -96 86599 -62 87575
rect 62 86599 96 87575
rect -34 86515 34 86549
rect -34 86407 34 86441
rect -96 85381 -62 86357
rect 62 85381 96 86357
rect -34 85297 34 85331
rect -34 85189 34 85223
rect -96 84163 -62 85139
rect 62 84163 96 85139
rect -34 84079 34 84113
rect -34 83971 34 84005
rect -96 82945 -62 83921
rect 62 82945 96 83921
rect -34 82861 34 82895
rect -34 82753 34 82787
rect -96 81727 -62 82703
rect 62 81727 96 82703
rect -34 81643 34 81677
rect -34 81535 34 81569
rect -96 80509 -62 81485
rect 62 80509 96 81485
rect -34 80425 34 80459
rect -34 80317 34 80351
rect -96 79291 -62 80267
rect 62 79291 96 80267
rect -34 79207 34 79241
rect -34 79099 34 79133
rect -96 78073 -62 79049
rect 62 78073 96 79049
rect -34 77989 34 78023
rect -34 77881 34 77915
rect -96 76855 -62 77831
rect 62 76855 96 77831
rect -34 76771 34 76805
rect -34 76663 34 76697
rect -96 75637 -62 76613
rect 62 75637 96 76613
rect -34 75553 34 75587
rect -34 75445 34 75479
rect -96 74419 -62 75395
rect 62 74419 96 75395
rect -34 74335 34 74369
rect -34 74227 34 74261
rect -96 73201 -62 74177
rect 62 73201 96 74177
rect -34 73117 34 73151
rect -34 73009 34 73043
rect -96 71983 -62 72959
rect 62 71983 96 72959
rect -34 71899 34 71933
rect -34 71791 34 71825
rect -96 70765 -62 71741
rect 62 70765 96 71741
rect -34 70681 34 70715
rect -34 70573 34 70607
rect -96 69547 -62 70523
rect 62 69547 96 70523
rect -34 69463 34 69497
rect -34 69355 34 69389
rect -96 68329 -62 69305
rect 62 68329 96 69305
rect -34 68245 34 68279
rect -34 68137 34 68171
rect -96 67111 -62 68087
rect 62 67111 96 68087
rect -34 67027 34 67061
rect -34 66919 34 66953
rect -96 65893 -62 66869
rect 62 65893 96 66869
rect -34 65809 34 65843
rect -34 65701 34 65735
rect -96 64675 -62 65651
rect 62 64675 96 65651
rect -34 64591 34 64625
rect -34 64483 34 64517
rect -96 63457 -62 64433
rect 62 63457 96 64433
rect -34 63373 34 63407
rect -34 63265 34 63299
rect -96 62239 -62 63215
rect 62 62239 96 63215
rect -34 62155 34 62189
rect -34 62047 34 62081
rect -96 61021 -62 61997
rect 62 61021 96 61997
rect -34 60937 34 60971
rect -34 60829 34 60863
rect -96 59803 -62 60779
rect 62 59803 96 60779
rect -34 59719 34 59753
rect -34 59611 34 59645
rect -96 58585 -62 59561
rect 62 58585 96 59561
rect -34 58501 34 58535
rect -34 58393 34 58427
rect -96 57367 -62 58343
rect 62 57367 96 58343
rect -34 57283 34 57317
rect -34 57175 34 57209
rect -96 56149 -62 57125
rect 62 56149 96 57125
rect -34 56065 34 56099
rect -34 55957 34 55991
rect -96 54931 -62 55907
rect 62 54931 96 55907
rect -34 54847 34 54881
rect -34 54739 34 54773
rect -96 53713 -62 54689
rect 62 53713 96 54689
rect -34 53629 34 53663
rect -34 53521 34 53555
rect -96 52495 -62 53471
rect 62 52495 96 53471
rect -34 52411 34 52445
rect -34 52303 34 52337
rect -96 51277 -62 52253
rect 62 51277 96 52253
rect -34 51193 34 51227
rect -34 51085 34 51119
rect -96 50059 -62 51035
rect 62 50059 96 51035
rect -34 49975 34 50009
rect -34 49867 34 49901
rect -96 48841 -62 49817
rect 62 48841 96 49817
rect -34 48757 34 48791
rect -34 48649 34 48683
rect -96 47623 -62 48599
rect 62 47623 96 48599
rect -34 47539 34 47573
rect -34 47431 34 47465
rect -96 46405 -62 47381
rect 62 46405 96 47381
rect -34 46321 34 46355
rect -34 46213 34 46247
rect -96 45187 -62 46163
rect 62 45187 96 46163
rect -34 45103 34 45137
rect -34 44995 34 45029
rect -96 43969 -62 44945
rect 62 43969 96 44945
rect -34 43885 34 43919
rect -34 43777 34 43811
rect -96 42751 -62 43727
rect 62 42751 96 43727
rect -34 42667 34 42701
rect -34 42559 34 42593
rect -96 41533 -62 42509
rect 62 41533 96 42509
rect -34 41449 34 41483
rect -34 41341 34 41375
rect -96 40315 -62 41291
rect 62 40315 96 41291
rect -34 40231 34 40265
rect -34 40123 34 40157
rect -96 39097 -62 40073
rect 62 39097 96 40073
rect -34 39013 34 39047
rect -34 38905 34 38939
rect -96 37879 -62 38855
rect 62 37879 96 38855
rect -34 37795 34 37829
rect -34 37687 34 37721
rect -96 36661 -62 37637
rect 62 36661 96 37637
rect -34 36577 34 36611
rect -34 36469 34 36503
rect -96 35443 -62 36419
rect 62 35443 96 36419
rect -34 35359 34 35393
rect -34 35251 34 35285
rect -96 34225 -62 35201
rect 62 34225 96 35201
rect -34 34141 34 34175
rect -34 34033 34 34067
rect -96 33007 -62 33983
rect 62 33007 96 33983
rect -34 32923 34 32957
rect -34 32815 34 32849
rect -96 31789 -62 32765
rect 62 31789 96 32765
rect -34 31705 34 31739
rect -34 31597 34 31631
rect -96 30571 -62 31547
rect 62 30571 96 31547
rect -34 30487 34 30521
rect -34 30379 34 30413
rect -96 29353 -62 30329
rect 62 29353 96 30329
rect -34 29269 34 29303
rect -34 29161 34 29195
rect -96 28135 -62 29111
rect 62 28135 96 29111
rect -34 28051 34 28085
rect -34 27943 34 27977
rect -96 26917 -62 27893
rect 62 26917 96 27893
rect -34 26833 34 26867
rect -34 26725 34 26759
rect -96 25699 -62 26675
rect 62 25699 96 26675
rect -34 25615 34 25649
rect -34 25507 34 25541
rect -96 24481 -62 25457
rect 62 24481 96 25457
rect -34 24397 34 24431
rect -34 24289 34 24323
rect -96 23263 -62 24239
rect 62 23263 96 24239
rect -34 23179 34 23213
rect -34 23071 34 23105
rect -96 22045 -62 23021
rect 62 22045 96 23021
rect -34 21961 34 21995
rect -34 21853 34 21887
rect -96 20827 -62 21803
rect 62 20827 96 21803
rect -34 20743 34 20777
rect -34 20635 34 20669
rect -96 19609 -62 20585
rect 62 19609 96 20585
rect -34 19525 34 19559
rect -34 19417 34 19451
rect -96 18391 -62 19367
rect 62 18391 96 19367
rect -34 18307 34 18341
rect -34 18199 34 18233
rect -96 17173 -62 18149
rect 62 17173 96 18149
rect -34 17089 34 17123
rect -34 16981 34 17015
rect -96 15955 -62 16931
rect 62 15955 96 16931
rect -34 15871 34 15905
rect -34 15763 34 15797
rect -96 14737 -62 15713
rect 62 14737 96 15713
rect -34 14653 34 14687
rect -34 14545 34 14579
rect -96 13519 -62 14495
rect 62 13519 96 14495
rect -34 13435 34 13469
rect -34 13327 34 13361
rect -96 12301 -62 13277
rect 62 12301 96 13277
rect -34 12217 34 12251
rect -34 12109 34 12143
rect -96 11083 -62 12059
rect 62 11083 96 12059
rect -34 10999 34 11033
rect -34 10891 34 10925
rect -96 9865 -62 10841
rect 62 9865 96 10841
rect -34 9781 34 9815
rect -34 9673 34 9707
rect -96 8647 -62 9623
rect 62 8647 96 9623
rect -34 8563 34 8597
rect -34 8455 34 8489
rect -96 7429 -62 8405
rect 62 7429 96 8405
rect -34 7345 34 7379
rect -34 7237 34 7271
rect -96 6211 -62 7187
rect 62 6211 96 7187
rect -34 6127 34 6161
rect -34 6019 34 6053
rect -96 4993 -62 5969
rect 62 4993 96 5969
rect -34 4909 34 4943
rect -34 4801 34 4835
rect -96 3775 -62 4751
rect 62 3775 96 4751
rect -34 3691 34 3725
rect -34 3583 34 3617
rect -96 2557 -62 3533
rect 62 2557 96 3533
rect -34 2473 34 2507
rect -34 2365 34 2399
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -96 121 -62 1097
rect 62 121 96 1097
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
rect -34 -2399 34 -2365
rect -34 -2507 34 -2473
rect -96 -3533 -62 -2557
rect 62 -3533 96 -2557
rect -34 -3617 34 -3583
rect -34 -3725 34 -3691
rect -96 -4751 -62 -3775
rect 62 -4751 96 -3775
rect -34 -4835 34 -4801
rect -34 -4943 34 -4909
rect -96 -5969 -62 -4993
rect 62 -5969 96 -4993
rect -34 -6053 34 -6019
rect -34 -6161 34 -6127
rect -96 -7187 -62 -6211
rect 62 -7187 96 -6211
rect -34 -7271 34 -7237
rect -34 -7379 34 -7345
rect -96 -8405 -62 -7429
rect 62 -8405 96 -7429
rect -34 -8489 34 -8455
rect -34 -8597 34 -8563
rect -96 -9623 -62 -8647
rect 62 -9623 96 -8647
rect -34 -9707 34 -9673
rect -34 -9815 34 -9781
rect -96 -10841 -62 -9865
rect 62 -10841 96 -9865
rect -34 -10925 34 -10891
rect -34 -11033 34 -10999
rect -96 -12059 -62 -11083
rect 62 -12059 96 -11083
rect -34 -12143 34 -12109
rect -34 -12251 34 -12217
rect -96 -13277 -62 -12301
rect 62 -13277 96 -12301
rect -34 -13361 34 -13327
rect -34 -13469 34 -13435
rect -96 -14495 -62 -13519
rect 62 -14495 96 -13519
rect -34 -14579 34 -14545
rect -34 -14687 34 -14653
rect -96 -15713 -62 -14737
rect 62 -15713 96 -14737
rect -34 -15797 34 -15763
rect -34 -15905 34 -15871
rect -96 -16931 -62 -15955
rect 62 -16931 96 -15955
rect -34 -17015 34 -16981
rect -34 -17123 34 -17089
rect -96 -18149 -62 -17173
rect 62 -18149 96 -17173
rect -34 -18233 34 -18199
rect -34 -18341 34 -18307
rect -96 -19367 -62 -18391
rect 62 -19367 96 -18391
rect -34 -19451 34 -19417
rect -34 -19559 34 -19525
rect -96 -20585 -62 -19609
rect 62 -20585 96 -19609
rect -34 -20669 34 -20635
rect -34 -20777 34 -20743
rect -96 -21803 -62 -20827
rect 62 -21803 96 -20827
rect -34 -21887 34 -21853
rect -34 -21995 34 -21961
rect -96 -23021 -62 -22045
rect 62 -23021 96 -22045
rect -34 -23105 34 -23071
rect -34 -23213 34 -23179
rect -96 -24239 -62 -23263
rect 62 -24239 96 -23263
rect -34 -24323 34 -24289
rect -34 -24431 34 -24397
rect -96 -25457 -62 -24481
rect 62 -25457 96 -24481
rect -34 -25541 34 -25507
rect -34 -25649 34 -25615
rect -96 -26675 -62 -25699
rect 62 -26675 96 -25699
rect -34 -26759 34 -26725
rect -34 -26867 34 -26833
rect -96 -27893 -62 -26917
rect 62 -27893 96 -26917
rect -34 -27977 34 -27943
rect -34 -28085 34 -28051
rect -96 -29111 -62 -28135
rect 62 -29111 96 -28135
rect -34 -29195 34 -29161
rect -34 -29303 34 -29269
rect -96 -30329 -62 -29353
rect 62 -30329 96 -29353
rect -34 -30413 34 -30379
rect -34 -30521 34 -30487
rect -96 -31547 -62 -30571
rect 62 -31547 96 -30571
rect -34 -31631 34 -31597
rect -34 -31739 34 -31705
rect -96 -32765 -62 -31789
rect 62 -32765 96 -31789
rect -34 -32849 34 -32815
rect -34 -32957 34 -32923
rect -96 -33983 -62 -33007
rect 62 -33983 96 -33007
rect -34 -34067 34 -34033
rect -34 -34175 34 -34141
rect -96 -35201 -62 -34225
rect 62 -35201 96 -34225
rect -34 -35285 34 -35251
rect -34 -35393 34 -35359
rect -96 -36419 -62 -35443
rect 62 -36419 96 -35443
rect -34 -36503 34 -36469
rect -34 -36611 34 -36577
rect -96 -37637 -62 -36661
rect 62 -37637 96 -36661
rect -34 -37721 34 -37687
rect -34 -37829 34 -37795
rect -96 -38855 -62 -37879
rect 62 -38855 96 -37879
rect -34 -38939 34 -38905
rect -34 -39047 34 -39013
rect -96 -40073 -62 -39097
rect 62 -40073 96 -39097
rect -34 -40157 34 -40123
rect -34 -40265 34 -40231
rect -96 -41291 -62 -40315
rect 62 -41291 96 -40315
rect -34 -41375 34 -41341
rect -34 -41483 34 -41449
rect -96 -42509 -62 -41533
rect 62 -42509 96 -41533
rect -34 -42593 34 -42559
rect -34 -42701 34 -42667
rect -96 -43727 -62 -42751
rect 62 -43727 96 -42751
rect -34 -43811 34 -43777
rect -34 -43919 34 -43885
rect -96 -44945 -62 -43969
rect 62 -44945 96 -43969
rect -34 -45029 34 -44995
rect -34 -45137 34 -45103
rect -96 -46163 -62 -45187
rect 62 -46163 96 -45187
rect -34 -46247 34 -46213
rect -34 -46355 34 -46321
rect -96 -47381 -62 -46405
rect 62 -47381 96 -46405
rect -34 -47465 34 -47431
rect -34 -47573 34 -47539
rect -96 -48599 -62 -47623
rect 62 -48599 96 -47623
rect -34 -48683 34 -48649
rect -34 -48791 34 -48757
rect -96 -49817 -62 -48841
rect 62 -49817 96 -48841
rect -34 -49901 34 -49867
rect -34 -50009 34 -49975
rect -96 -51035 -62 -50059
rect 62 -51035 96 -50059
rect -34 -51119 34 -51085
rect -34 -51227 34 -51193
rect -96 -52253 -62 -51277
rect 62 -52253 96 -51277
rect -34 -52337 34 -52303
rect -34 -52445 34 -52411
rect -96 -53471 -62 -52495
rect 62 -53471 96 -52495
rect -34 -53555 34 -53521
rect -34 -53663 34 -53629
rect -96 -54689 -62 -53713
rect 62 -54689 96 -53713
rect -34 -54773 34 -54739
rect -34 -54881 34 -54847
rect -96 -55907 -62 -54931
rect 62 -55907 96 -54931
rect -34 -55991 34 -55957
rect -34 -56099 34 -56065
rect -96 -57125 -62 -56149
rect 62 -57125 96 -56149
rect -34 -57209 34 -57175
rect -34 -57317 34 -57283
rect -96 -58343 -62 -57367
rect 62 -58343 96 -57367
rect -34 -58427 34 -58393
rect -34 -58535 34 -58501
rect -96 -59561 -62 -58585
rect 62 -59561 96 -58585
rect -34 -59645 34 -59611
rect -34 -59753 34 -59719
rect -96 -60779 -62 -59803
rect 62 -60779 96 -59803
rect -34 -60863 34 -60829
rect -34 -60971 34 -60937
rect -96 -61997 -62 -61021
rect 62 -61997 96 -61021
rect -34 -62081 34 -62047
rect -34 -62189 34 -62155
rect -96 -63215 -62 -62239
rect 62 -63215 96 -62239
rect -34 -63299 34 -63265
rect -34 -63407 34 -63373
rect -96 -64433 -62 -63457
rect 62 -64433 96 -63457
rect -34 -64517 34 -64483
rect -34 -64625 34 -64591
rect -96 -65651 -62 -64675
rect 62 -65651 96 -64675
rect -34 -65735 34 -65701
rect -34 -65843 34 -65809
rect -96 -66869 -62 -65893
rect 62 -66869 96 -65893
rect -34 -66953 34 -66919
rect -34 -67061 34 -67027
rect -96 -68087 -62 -67111
rect 62 -68087 96 -67111
rect -34 -68171 34 -68137
rect -34 -68279 34 -68245
rect -96 -69305 -62 -68329
rect 62 -69305 96 -68329
rect -34 -69389 34 -69355
rect -34 -69497 34 -69463
rect -96 -70523 -62 -69547
rect 62 -70523 96 -69547
rect -34 -70607 34 -70573
rect -34 -70715 34 -70681
rect -96 -71741 -62 -70765
rect 62 -71741 96 -70765
rect -34 -71825 34 -71791
rect -34 -71933 34 -71899
rect -96 -72959 -62 -71983
rect 62 -72959 96 -71983
rect -34 -73043 34 -73009
rect -34 -73151 34 -73117
rect -96 -74177 -62 -73201
rect 62 -74177 96 -73201
rect -34 -74261 34 -74227
rect -34 -74369 34 -74335
rect -96 -75395 -62 -74419
rect 62 -75395 96 -74419
rect -34 -75479 34 -75445
rect -34 -75587 34 -75553
rect -96 -76613 -62 -75637
rect 62 -76613 96 -75637
rect -34 -76697 34 -76663
rect -34 -76805 34 -76771
rect -96 -77831 -62 -76855
rect 62 -77831 96 -76855
rect -34 -77915 34 -77881
rect -34 -78023 34 -77989
rect -96 -79049 -62 -78073
rect 62 -79049 96 -78073
rect -34 -79133 34 -79099
rect -34 -79241 34 -79207
rect -96 -80267 -62 -79291
rect 62 -80267 96 -79291
rect -34 -80351 34 -80317
rect -34 -80459 34 -80425
rect -96 -81485 -62 -80509
rect 62 -81485 96 -80509
rect -34 -81569 34 -81535
rect -34 -81677 34 -81643
rect -96 -82703 -62 -81727
rect 62 -82703 96 -81727
rect -34 -82787 34 -82753
rect -34 -82895 34 -82861
rect -96 -83921 -62 -82945
rect 62 -83921 96 -82945
rect -34 -84005 34 -83971
rect -34 -84113 34 -84079
rect -96 -85139 -62 -84163
rect 62 -85139 96 -84163
rect -34 -85223 34 -85189
rect -34 -85331 34 -85297
rect -96 -86357 -62 -85381
rect 62 -86357 96 -85381
rect -34 -86441 34 -86407
rect -34 -86549 34 -86515
rect -96 -87575 -62 -86599
rect 62 -87575 96 -86599
rect -34 -87659 34 -87625
rect -34 -87767 34 -87733
rect -96 -88793 -62 -87817
rect 62 -88793 96 -87817
rect -34 -88877 34 -88843
rect -34 -88985 34 -88951
rect -96 -90011 -62 -89035
rect 62 -90011 96 -89035
rect -34 -90095 34 -90061
rect -34 -90203 34 -90169
rect -96 -91229 -62 -90253
rect 62 -91229 96 -90253
rect -34 -91313 34 -91279
rect -34 -91421 34 -91387
rect -96 -92447 -62 -91471
rect 62 -92447 96 -91471
rect -34 -92531 34 -92497
rect -34 -92639 34 -92605
rect -96 -93665 -62 -92689
rect 62 -93665 96 -92689
rect -34 -93749 34 -93715
rect -34 -93857 34 -93823
rect -96 -94883 -62 -93907
rect 62 -94883 96 -93907
rect -34 -94967 34 -94933
rect -34 -95075 34 -95041
rect -96 -96101 -62 -95125
rect 62 -96101 96 -95125
rect -34 -96185 34 -96151
rect -34 -96293 34 -96259
rect -96 -97319 -62 -96343
rect 62 -97319 96 -96343
rect -34 -97403 34 -97369
rect -34 -97511 34 -97477
rect -96 -98537 -62 -97561
rect 62 -98537 96 -97561
rect -34 -98621 34 -98587
rect -34 -98729 34 -98695
rect -96 -99755 -62 -98779
rect 62 -99755 96 -98779
rect -34 -99839 34 -99805
rect -34 -99947 34 -99913
rect -96 -100973 -62 -99997
rect 62 -100973 96 -99997
rect -34 -101057 34 -101023
rect -34 -101165 34 -101131
rect -96 -102191 -62 -101215
rect 62 -102191 96 -101215
rect -34 -102275 34 -102241
rect -34 -102383 34 -102349
rect -96 -103409 -62 -102433
rect 62 -103409 96 -102433
rect -34 -103493 34 -103459
rect -34 -103601 34 -103567
rect -96 -104627 -62 -103651
rect 62 -104627 96 -103651
rect -34 -104711 34 -104677
rect -34 -104819 34 -104785
rect -96 -105845 -62 -104869
rect 62 -105845 96 -104869
rect -34 -105929 34 -105895
rect -34 -106037 34 -106003
rect -96 -107063 -62 -106087
rect 62 -107063 96 -106087
rect -34 -107147 34 -107113
rect -34 -107255 34 -107221
rect -96 -108281 -62 -107305
rect 62 -108281 96 -107305
rect -34 -108365 34 -108331
rect -34 -108473 34 -108439
rect -96 -109499 -62 -108523
rect 62 -109499 96 -108523
rect -34 -109583 34 -109549
rect -34 -109691 34 -109657
rect -96 -110717 -62 -109741
rect 62 -110717 96 -109741
rect -34 -110801 34 -110767
rect -34 -110909 34 -110875
rect -96 -111935 -62 -110959
rect 62 -111935 96 -110959
rect -34 -112019 34 -111985
rect -34 -112127 34 -112093
rect -96 -113153 -62 -112177
rect 62 -113153 96 -112177
rect -34 -113237 34 -113203
rect -34 -113345 34 -113311
rect -96 -114371 -62 -113395
rect 62 -114371 96 -113395
rect -34 -114455 34 -114421
rect -34 -114563 34 -114529
rect -96 -115589 -62 -114613
rect 62 -115589 96 -114613
rect -34 -115673 34 -115639
rect -34 -115781 34 -115747
rect -96 -116807 -62 -115831
rect 62 -116807 96 -115831
rect -34 -116891 34 -116857
rect -34 -116999 34 -116965
rect -96 -118025 -62 -117049
rect 62 -118025 96 -117049
rect -34 -118109 34 -118075
rect -34 -118217 34 -118183
rect -96 -119243 -62 -118267
rect 62 -119243 96 -118267
rect -34 -119327 34 -119293
rect -34 -119435 34 -119401
rect -96 -120461 -62 -119485
rect 62 -120461 96 -119485
rect -34 -120545 34 -120511
rect -34 -120653 34 -120619
rect -96 -121679 -62 -120703
rect 62 -121679 96 -120703
rect -34 -121763 34 -121729
rect -34 -121871 34 -121837
rect -96 -122897 -62 -121921
rect 62 -122897 96 -121921
rect -34 -122981 34 -122947
rect -34 -123089 34 -123055
rect -96 -124115 -62 -123139
rect 62 -124115 96 -123139
rect -34 -124199 34 -124165
rect -34 -124307 34 -124273
rect -96 -125333 -62 -124357
rect 62 -125333 96 -124357
rect -34 -125417 34 -125383
rect -34 -125525 34 -125491
rect -96 -126551 -62 -125575
rect 62 -126551 96 -125575
rect -34 -126635 34 -126601
rect -34 -126743 34 -126709
rect -96 -127769 -62 -126793
rect 62 -127769 96 -126793
rect -34 -127853 34 -127819
rect -34 -127961 34 -127927
rect -96 -128987 -62 -128011
rect 62 -128987 96 -128011
rect -34 -129071 34 -129037
rect -34 -129179 34 -129145
rect -96 -130205 -62 -129229
rect 62 -130205 96 -129229
rect -34 -130289 34 -130255
rect -34 -130397 34 -130363
rect -96 -131423 -62 -130447
rect 62 -131423 96 -130447
rect -34 -131507 34 -131473
rect -34 -131615 34 -131581
rect -96 -132641 -62 -131665
rect 62 -132641 96 -131665
rect -34 -132725 34 -132691
rect -34 -132833 34 -132799
rect -96 -133859 -62 -132883
rect 62 -133859 96 -132883
rect -34 -133943 34 -133909
rect -34 -134051 34 -134017
rect -96 -135077 -62 -134101
rect 62 -135077 96 -134101
rect -34 -135161 34 -135127
rect -34 -135269 34 -135235
rect -96 -136295 -62 -135319
rect 62 -136295 96 -135319
rect -34 -136379 34 -136345
rect -34 -136487 34 -136453
rect -96 -137513 -62 -136537
rect 62 -137513 96 -136537
rect -34 -137597 34 -137563
rect -34 -137705 34 -137671
rect -96 -138731 -62 -137755
rect 62 -138731 96 -137755
rect -34 -138815 34 -138781
rect -34 -138923 34 -138889
rect -96 -139949 -62 -138973
rect 62 -139949 96 -138973
rect -34 -140033 34 -139999
rect -34 -140141 34 -140107
rect -96 -141167 -62 -140191
rect 62 -141167 96 -140191
rect -34 -141251 34 -141217
rect -34 -141359 34 -141325
rect -96 -142385 -62 -141409
rect 62 -142385 96 -141409
rect -34 -142469 34 -142435
rect -34 -142577 34 -142543
rect -96 -143603 -62 -142627
rect 62 -143603 96 -142627
rect -34 -143687 34 -143653
rect -34 -143795 34 -143761
rect -96 -144821 -62 -143845
rect 62 -144821 96 -143845
rect -34 -144905 34 -144871
rect -34 -145013 34 -144979
rect -96 -146039 -62 -145063
rect 62 -146039 96 -145063
rect -34 -146123 34 -146089
rect -34 -146231 34 -146197
rect -96 -147257 -62 -146281
rect 62 -147257 96 -146281
rect -34 -147341 34 -147307
rect -34 -147449 34 -147415
rect -96 -148475 -62 -147499
rect 62 -148475 96 -147499
rect -34 -148559 34 -148525
rect -34 -148667 34 -148633
rect -96 -149693 -62 -148717
rect 62 -149693 96 -148717
rect -34 -149777 34 -149743
rect -34 -149885 34 -149851
rect -96 -150911 -62 -149935
rect 62 -150911 96 -149935
rect -34 -150995 34 -150961
rect -34 -151103 34 -151069
rect -96 -152129 -62 -151153
rect 62 -152129 96 -151153
rect -34 -152213 34 -152179
rect -34 -152321 34 -152287
rect -96 -153347 -62 -152371
rect 62 -153347 96 -152371
rect -34 -153431 34 -153397
rect -34 -153539 34 -153505
rect -96 -154565 -62 -153589
rect 62 -154565 96 -153589
rect -34 -154649 34 -154615
rect -34 -154757 34 -154723
rect -96 -155783 -62 -154807
rect 62 -155783 96 -154807
rect -34 -155867 34 -155833
rect -34 -155975 34 -155941
rect -96 -157001 -62 -156025
rect 62 -157001 96 -156025
rect -34 -157085 34 -157051
rect -34 -157193 34 -157159
rect -96 -158219 -62 -157243
rect 62 -158219 96 -157243
rect -34 -158303 34 -158269
rect -34 -158411 34 -158377
rect -96 -159437 -62 -158461
rect 62 -159437 96 -158461
rect -34 -159521 34 -159487
rect -34 -159629 34 -159595
rect -96 -160655 -62 -159679
rect 62 -160655 96 -159679
rect -34 -160739 34 -160705
rect -34 -160847 34 -160813
rect -96 -161873 -62 -160897
rect 62 -161873 96 -160897
rect -34 -161957 34 -161923
rect -34 -162065 34 -162031
rect -96 -163091 -62 -162115
rect 62 -163091 96 -162115
rect -34 -163175 34 -163141
rect -34 -163283 34 -163249
rect -96 -164309 -62 -163333
rect 62 -164309 96 -163333
rect -34 -164393 34 -164359
rect -34 -164501 34 -164467
rect -96 -165527 -62 -164551
rect 62 -165527 96 -164551
rect -34 -165611 34 -165577
rect -34 -165719 34 -165685
rect -96 -166745 -62 -165769
rect 62 -166745 96 -165769
rect -34 -166829 34 -166795
rect -34 -166937 34 -166903
rect -96 -167963 -62 -166987
rect 62 -167963 96 -166987
rect -34 -168047 34 -168013
rect -34 -168155 34 -168121
rect -96 -169181 -62 -168205
rect 62 -169181 96 -168205
rect -34 -169265 34 -169231
rect -34 -169373 34 -169339
rect -96 -170399 -62 -169423
rect 62 -170399 96 -169423
rect -34 -170483 34 -170449
rect -34 -170591 34 -170557
rect -96 -171617 -62 -170641
rect 62 -171617 96 -170641
rect -34 -171701 34 -171667
rect -34 -171809 34 -171775
rect -96 -172835 -62 -171859
rect 62 -172835 96 -171859
rect -34 -172919 34 -172885
rect -34 -173027 34 -172993
rect -96 -174053 -62 -173077
rect 62 -174053 96 -173077
rect -34 -174137 34 -174103
rect -34 -174245 34 -174211
rect -96 -175271 -62 -174295
rect 62 -175271 96 -174295
rect -34 -175355 34 -175321
rect -34 -175463 34 -175429
rect -96 -176489 -62 -175513
rect 62 -176489 96 -175513
rect -34 -176573 34 -176539
rect -34 -176681 34 -176647
rect -96 -177707 -62 -176731
rect 62 -177707 96 -176731
rect -34 -177791 34 -177757
rect -34 -177899 34 -177865
rect -96 -178925 -62 -177949
rect 62 -178925 96 -177949
rect -34 -179009 34 -178975
rect -34 -179117 34 -179083
rect -96 -180143 -62 -179167
rect 62 -180143 96 -179167
rect -34 -180227 34 -180193
rect -34 -180335 34 -180301
rect -96 -181361 -62 -180385
rect 62 -181361 96 -180385
rect -34 -181445 34 -181411
rect -34 -181553 34 -181519
rect -96 -182579 -62 -181603
rect 62 -182579 96 -181603
rect -34 -182663 34 -182629
rect -34 -182771 34 -182737
rect -96 -183797 -62 -182821
rect 62 -183797 96 -182821
rect -34 -183881 34 -183847
rect -34 -183989 34 -183955
rect -96 -185015 -62 -184039
rect 62 -185015 96 -184039
rect -34 -185099 34 -185065
rect -34 -185207 34 -185173
rect -96 -186233 -62 -185257
rect 62 -186233 96 -185257
rect -34 -186317 34 -186283
rect -34 -186425 34 -186391
rect -96 -187451 -62 -186475
rect 62 -187451 96 -186475
rect -34 -187535 34 -187501
rect -34 -187643 34 -187609
rect -96 -188669 -62 -187693
rect 62 -188669 96 -187693
rect -34 -188753 34 -188719
rect -34 -188861 34 -188827
rect -96 -189887 -62 -188911
rect 62 -189887 96 -188911
rect -34 -189971 34 -189937
rect -34 -190079 34 -190045
rect -96 -191105 -62 -190129
rect 62 -191105 96 -190129
rect -34 -191189 34 -191155
rect -34 -191297 34 -191263
rect -96 -192323 -62 -191347
rect 62 -192323 96 -191347
rect -34 -192407 34 -192373
rect -34 -192515 34 -192481
rect -96 -193541 -62 -192565
rect 62 -193541 96 -192565
rect -34 -193625 34 -193591
rect -34 -193733 34 -193699
rect -96 -194759 -62 -193783
rect 62 -194759 96 -193783
rect -34 -194843 34 -194809
rect -34 -194951 34 -194917
rect -96 -195977 -62 -195001
rect 62 -195977 96 -195001
rect -34 -196061 34 -196027
rect -34 -196169 34 -196135
rect -96 -197195 -62 -196219
rect 62 -197195 96 -196219
rect -34 -197279 34 -197245
rect -34 -197387 34 -197353
rect -96 -198413 -62 -197437
rect 62 -198413 96 -197437
rect -34 -198497 34 -198463
rect -34 -198605 34 -198571
rect -96 -199631 -62 -198655
rect 62 -199631 96 -198655
rect -34 -199715 34 -199681
rect -34 -199823 34 -199789
rect -96 -200849 -62 -199873
rect 62 -200849 96 -199873
rect -34 -200933 34 -200899
rect -34 -201041 34 -201007
rect -96 -202067 -62 -201091
rect 62 -202067 96 -201091
rect -34 -202151 34 -202117
rect -34 -202259 34 -202225
rect -96 -203285 -62 -202309
rect 62 -203285 96 -202309
rect -34 -203369 34 -203335
rect -34 -203477 34 -203443
rect -96 -204503 -62 -203527
rect 62 -204503 96 -203527
rect -34 -204587 34 -204553
rect -34 -204695 34 -204661
rect -96 -205721 -62 -204745
rect 62 -205721 96 -204745
rect -34 -205805 34 -205771
rect -34 -205913 34 -205879
rect -96 -206939 -62 -205963
rect 62 -206939 96 -205963
rect -34 -207023 34 -206989
rect -34 -207131 34 -207097
rect -96 -208157 -62 -207181
rect 62 -208157 96 -207181
rect -34 -208241 34 -208207
rect -34 -208349 34 -208315
rect -96 -209375 -62 -208399
rect 62 -209375 96 -208399
rect -34 -209459 34 -209425
rect -34 -209567 34 -209533
rect -96 -210593 -62 -209617
rect 62 -210593 96 -209617
rect -34 -210677 34 -210643
rect -34 -210785 34 -210751
rect -96 -211811 -62 -210835
rect 62 -211811 96 -210835
rect -34 -211895 34 -211861
rect -34 -212003 34 -211969
rect -96 -213029 -62 -212053
rect 62 -213029 96 -212053
rect -34 -213113 34 -213079
rect -34 -213221 34 -213187
rect -96 -214247 -62 -213271
rect 62 -214247 96 -213271
rect -34 -214331 34 -214297
rect -34 -214439 34 -214405
rect -96 -215465 -62 -214489
rect 62 -215465 96 -214489
rect -34 -215549 34 -215515
rect -34 -215657 34 -215623
rect -96 -216683 -62 -215707
rect 62 -216683 96 -215707
rect -34 -216767 34 -216733
rect -34 -216875 34 -216841
rect -96 -217901 -62 -216925
rect 62 -217901 96 -216925
rect -34 -217985 34 -217951
rect -34 -218093 34 -218059
rect -96 -219119 -62 -218143
rect 62 -219119 96 -218143
rect -34 -219203 34 -219169
rect -34 -219311 34 -219277
rect -96 -220337 -62 -219361
rect 62 -220337 96 -219361
rect -34 -220421 34 -220387
rect -34 -220529 34 -220495
rect -96 -221555 -62 -220579
rect 62 -221555 96 -220579
rect -34 -221639 34 -221605
rect -34 -221747 34 -221713
rect -96 -222773 -62 -221797
rect 62 -222773 96 -221797
rect -34 -222857 34 -222823
rect -34 -222965 34 -222931
rect -96 -223991 -62 -223015
rect 62 -223991 96 -223015
rect -34 -224075 34 -224041
rect -34 -224183 34 -224149
rect -96 -225209 -62 -224233
rect 62 -225209 96 -224233
rect -34 -225293 34 -225259
rect -34 -225401 34 -225367
rect -96 -226427 -62 -225451
rect 62 -226427 96 -225451
rect -34 -226511 34 -226477
rect -34 -226619 34 -226585
rect -96 -227645 -62 -226669
rect 62 -227645 96 -226669
rect -34 -227729 34 -227695
rect -34 -227837 34 -227803
rect -96 -228863 -62 -227887
rect 62 -228863 96 -227887
rect -34 -228947 34 -228913
rect -34 -229055 34 -229021
rect -96 -230081 -62 -229105
rect 62 -230081 96 -229105
rect -34 -230165 34 -230131
rect -34 -230273 34 -230239
rect -96 -231299 -62 -230323
rect 62 -231299 96 -230323
rect -34 -231383 34 -231349
rect -34 -231491 34 -231457
rect -96 -232517 -62 -231541
rect 62 -232517 96 -231541
rect -34 -232601 34 -232567
rect -34 -232709 34 -232675
rect -96 -233735 -62 -232759
rect 62 -233735 96 -232759
rect -34 -233819 34 -233785
rect -34 -233927 34 -233893
rect -96 -234953 -62 -233977
rect 62 -234953 96 -233977
rect -34 -235037 34 -235003
rect -34 -235145 34 -235111
rect -96 -236171 -62 -235195
rect 62 -236171 96 -235195
rect -34 -236255 34 -236221
rect -34 -236363 34 -236329
rect -96 -237389 -62 -236413
rect 62 -237389 96 -236413
rect -34 -237473 34 -237439
rect -34 -237581 34 -237547
rect -96 -238607 -62 -237631
rect 62 -238607 96 -237631
rect -34 -238691 34 -238657
rect -34 -238799 34 -238765
rect -96 -239825 -62 -238849
rect 62 -239825 96 -238849
rect -34 -239909 34 -239875
rect -34 -240017 34 -239983
rect -96 -241043 -62 -240067
rect 62 -241043 96 -240067
rect -34 -241127 34 -241093
rect -34 -241235 34 -241201
rect -96 -242261 -62 -241285
rect 62 -242261 96 -241285
rect -34 -242345 34 -242311
rect -34 -242453 34 -242419
rect -96 -243479 -62 -242503
rect 62 -243479 96 -242503
rect -34 -243563 34 -243529
rect -34 -243671 34 -243637
rect -96 -244697 -62 -243721
rect 62 -244697 96 -243721
rect -34 -244781 34 -244747
rect -34 -244889 34 -244855
rect -96 -245915 -62 -244939
rect 62 -245915 96 -244939
rect -34 -245999 34 -245965
rect -34 -246107 34 -246073
rect -96 -247133 -62 -246157
rect 62 -247133 96 -246157
rect -34 -247217 34 -247183
rect -34 -247325 34 -247291
rect -96 -248351 -62 -247375
rect 62 -248351 96 -247375
rect -34 -248435 34 -248401
rect -34 -248543 34 -248509
rect -96 -249569 -62 -248593
rect 62 -249569 96 -248593
rect -34 -249653 34 -249619
rect -34 -249761 34 -249727
rect -96 -250787 -62 -249811
rect 62 -250787 96 -249811
rect -34 -250871 34 -250837
rect -34 -250979 34 -250945
rect -96 -252005 -62 -251029
rect 62 -252005 96 -251029
rect -34 -252089 34 -252055
rect -34 -252197 34 -252163
rect -96 -253223 -62 -252247
rect 62 -253223 96 -252247
rect -34 -253307 34 -253273
rect -34 -253415 34 -253381
rect -96 -254441 -62 -253465
rect 62 -254441 96 -253465
rect -34 -254525 34 -254491
rect -34 -254633 34 -254599
rect -96 -255659 -62 -254683
rect 62 -255659 96 -254683
rect -34 -255743 34 -255709
rect -34 -255851 34 -255817
rect -96 -256877 -62 -255901
rect 62 -256877 96 -255901
rect -34 -256961 34 -256927
rect -34 -257069 34 -257035
rect -96 -258095 -62 -257119
rect 62 -258095 96 -257119
rect -34 -258179 34 -258145
rect -34 -258287 34 -258253
rect -96 -259313 -62 -258337
rect 62 -259313 96 -258337
rect -34 -259397 34 -259363
rect -34 -259505 34 -259471
rect -96 -260531 -62 -259555
rect 62 -260531 96 -259555
rect -34 -260615 34 -260581
rect -34 -260723 34 -260689
rect -96 -261749 -62 -260773
rect 62 -261749 96 -260773
rect -34 -261833 34 -261799
rect -34 -261941 34 -261907
rect -96 -262967 -62 -261991
rect 62 -262967 96 -261991
rect -34 -263051 34 -263017
rect -34 -263159 34 -263125
rect -96 -264185 -62 -263209
rect 62 -264185 96 -263209
rect -34 -264269 34 -264235
rect -34 -264377 34 -264343
rect -96 -265403 -62 -264427
rect 62 -265403 96 -264427
rect -34 -265487 34 -265453
rect -34 -265595 34 -265561
rect -96 -266621 -62 -265645
rect 62 -266621 96 -265645
rect -34 -266705 34 -266671
rect -34 -266813 34 -266779
rect -96 -267839 -62 -266863
rect 62 -267839 96 -266863
rect -34 -267923 34 -267889
rect -34 -268031 34 -267997
rect -96 -269057 -62 -268081
rect 62 -269057 96 -268081
rect -34 -269141 34 -269107
rect -34 -269249 34 -269215
rect -96 -270275 -62 -269299
rect 62 -270275 96 -269299
rect -34 -270359 34 -270325
rect -34 -270467 34 -270433
rect -96 -271493 -62 -270517
rect 62 -271493 96 -270517
rect -34 -271577 34 -271543
rect -34 -271685 34 -271651
rect -96 -272711 -62 -271735
rect 62 -272711 96 -271735
rect -34 -272795 34 -272761
rect -34 -272903 34 -272869
rect -96 -273929 -62 -272953
rect 62 -273929 96 -272953
rect -34 -274013 34 -273979
rect -34 -274121 34 -274087
rect -96 -275147 -62 -274171
rect 62 -275147 96 -274171
rect -34 -275231 34 -275197
rect -34 -275339 34 -275305
rect -96 -276365 -62 -275389
rect 62 -276365 96 -275389
rect -34 -276449 34 -276415
rect -34 -276557 34 -276523
rect -96 -277583 -62 -276607
rect 62 -277583 96 -276607
rect -34 -277667 34 -277633
rect -34 -277775 34 -277741
rect -96 -278801 -62 -277825
rect 62 -278801 96 -277825
rect -34 -278885 34 -278851
rect -34 -278993 34 -278959
rect -96 -280019 -62 -279043
rect 62 -280019 96 -279043
rect -34 -280103 34 -280069
rect -34 -280211 34 -280177
rect -96 -281237 -62 -280261
rect 62 -281237 96 -280261
rect -34 -281321 34 -281287
rect -34 -281429 34 -281395
rect -96 -282455 -62 -281479
rect 62 -282455 96 -281479
rect -34 -282539 34 -282505
rect -34 -282647 34 -282613
rect -96 -283673 -62 -282697
rect 62 -283673 96 -282697
rect -34 -283757 34 -283723
rect -34 -283865 34 -283831
rect -96 -284891 -62 -283915
rect 62 -284891 96 -283915
rect -34 -284975 34 -284941
rect -34 -285083 34 -285049
rect -96 -286109 -62 -285133
rect 62 -286109 96 -285133
rect -34 -286193 34 -286159
rect -34 -286301 34 -286267
rect -96 -287327 -62 -286351
rect 62 -287327 96 -286351
rect -34 -287411 34 -287377
rect -34 -287519 34 -287485
rect -96 -288545 -62 -287569
rect 62 -288545 96 -287569
rect -34 -288629 34 -288595
rect -34 -288737 34 -288703
rect -96 -289763 -62 -288787
rect 62 -289763 96 -288787
rect -34 -289847 34 -289813
rect -34 -289955 34 -289921
rect -96 -290981 -62 -290005
rect 62 -290981 96 -290005
rect -34 -291065 34 -291031
rect -34 -291173 34 -291139
rect -96 -292199 -62 -291223
rect 62 -292199 96 -291223
rect -34 -292283 34 -292249
rect -34 -292391 34 -292357
rect -96 -293417 -62 -292441
rect 62 -293417 96 -292441
rect -34 -293501 34 -293467
rect -34 -293609 34 -293575
rect -96 -294635 -62 -293659
rect 62 -294635 96 -293659
rect -34 -294719 34 -294685
rect -34 -294827 34 -294793
rect -96 -295853 -62 -294877
rect 62 -295853 96 -294877
rect -34 -295937 34 -295903
rect -34 -296045 34 -296011
rect -96 -297071 -62 -296095
rect 62 -297071 96 -296095
rect -34 -297155 34 -297121
rect -34 -297263 34 -297229
rect -96 -298289 -62 -297313
rect 62 -298289 96 -297313
rect -34 -298373 34 -298339
rect -34 -298481 34 -298447
rect -96 -299507 -62 -298531
rect 62 -299507 96 -298531
rect -34 -299591 34 -299557
rect -34 -299699 34 -299665
rect -96 -300725 -62 -299749
rect 62 -300725 96 -299749
rect -34 -300809 34 -300775
rect -34 -300917 34 -300883
rect -96 -301943 -62 -300967
rect 62 -301943 96 -300967
rect -34 -302027 34 -301993
rect -34 -302135 34 -302101
rect -96 -303161 -62 -302185
rect 62 -303161 96 -302185
rect -34 -303245 34 -303211
rect -34 -303353 34 -303319
rect -96 -304379 -62 -303403
rect 62 -304379 96 -303403
rect -34 -304463 34 -304429
rect -34 -304571 34 -304537
rect -96 -305597 -62 -304621
rect 62 -305597 96 -304621
rect -34 -305681 34 -305647
rect -34 -305789 34 -305755
rect -96 -306815 -62 -305839
rect 62 -306815 96 -305839
rect -34 -306899 34 -306865
rect -34 -307007 34 -306973
rect -96 -308033 -62 -307057
rect 62 -308033 96 -307057
rect -34 -308117 34 -308083
rect -34 -308225 34 -308191
rect -96 -309251 -62 -308275
rect 62 -309251 96 -308275
rect -34 -309335 34 -309301
rect -34 -309443 34 -309409
rect -96 -310469 -62 -309493
rect 62 -310469 96 -309493
rect -34 -310553 34 -310519
rect -34 -310661 34 -310627
rect -96 -311687 -62 -310711
rect 62 -311687 96 -310711
rect -34 -311771 34 -311737
rect -34 -311879 34 -311845
rect -96 -312905 -62 -311929
rect 62 -312905 96 -311929
rect -34 -312989 34 -312955
rect -34 -313097 34 -313063
rect -96 -314123 -62 -313147
rect 62 -314123 96 -313147
rect -34 -314207 34 -314173
rect -34 -314315 34 -314281
rect -96 -315341 -62 -314365
rect 62 -315341 96 -314365
rect -34 -315425 34 -315391
rect -34 -315533 34 -315499
rect -96 -316559 -62 -315583
rect 62 -316559 96 -315583
rect -34 -316643 34 -316609
rect -34 -316751 34 -316717
rect -96 -317777 -62 -316801
rect 62 -317777 96 -316801
rect -34 -317861 34 -317827
rect -34 -317969 34 -317935
rect -96 -318995 -62 -318019
rect 62 -318995 96 -318019
rect -34 -319079 34 -319045
rect -34 -319187 34 -319153
rect -96 -320213 -62 -319237
rect 62 -320213 96 -319237
rect -34 -320297 34 -320263
rect -34 -320405 34 -320371
rect -96 -321431 -62 -320455
rect 62 -321431 96 -320455
rect -34 -321515 34 -321481
rect -34 -321623 34 -321589
rect -96 -322649 -62 -321673
rect 62 -322649 96 -321673
rect -34 -322733 34 -322699
rect -34 -322841 34 -322807
rect -96 -323867 -62 -322891
rect 62 -323867 96 -322891
rect -34 -323951 34 -323917
rect -34 -324059 34 -324025
rect -96 -325085 -62 -324109
rect 62 -325085 96 -324109
rect -34 -325169 34 -325135
rect -34 -325277 34 -325243
rect -96 -326303 -62 -325327
rect 62 -326303 96 -325327
rect -34 -326387 34 -326353
rect -34 -326495 34 -326461
rect -96 -327521 -62 -326545
rect 62 -327521 96 -326545
rect -34 -327605 34 -327571
rect -34 -327713 34 -327679
rect -96 -328739 -62 -327763
rect 62 -328739 96 -327763
rect -34 -328823 34 -328789
rect -34 -328931 34 -328897
rect -96 -329957 -62 -328981
rect 62 -329957 96 -328981
rect -34 -330041 34 -330007
rect -34 -330149 34 -330115
rect -96 -331175 -62 -330199
rect 62 -331175 96 -330199
rect -34 -331259 34 -331225
rect -34 -331367 34 -331333
rect -96 -332393 -62 -331417
rect 62 -332393 96 -331417
rect -34 -332477 34 -332443
rect -34 -332585 34 -332551
rect -96 -333611 -62 -332635
rect 62 -333611 96 -332635
rect -34 -333695 34 -333661
rect -34 -333803 34 -333769
rect -96 -334829 -62 -333853
rect 62 -334829 96 -333853
rect -34 -334913 34 -334879
rect -34 -335021 34 -334987
rect -96 -336047 -62 -335071
rect 62 -336047 96 -335071
rect -34 -336131 34 -336097
rect -34 -336239 34 -336205
rect -96 -337265 -62 -336289
rect 62 -337265 96 -336289
rect -34 -337349 34 -337315
rect -34 -337457 34 -337423
rect -96 -338483 -62 -337507
rect 62 -338483 96 -337507
rect -34 -338567 34 -338533
rect -34 -338675 34 -338641
rect -96 -339701 -62 -338725
rect 62 -339701 96 -338725
rect -34 -339785 34 -339751
rect -34 -339893 34 -339859
rect -96 -340919 -62 -339943
rect 62 -340919 96 -339943
rect -34 -341003 34 -340969
rect -34 -341111 34 -341077
rect -96 -342137 -62 -341161
rect 62 -342137 96 -341161
rect -34 -342221 34 -342187
rect -34 -342329 34 -342295
rect -96 -343355 -62 -342379
rect 62 -343355 96 -342379
rect -34 -343439 34 -343405
rect -34 -343547 34 -343513
rect -96 -344573 -62 -343597
rect 62 -344573 96 -343597
rect -34 -344657 34 -344623
rect -34 -344765 34 -344731
rect -96 -345791 -62 -344815
rect 62 -345791 96 -344815
rect -34 -345875 34 -345841
rect -34 -345983 34 -345949
rect -96 -347009 -62 -346033
rect 62 -347009 96 -346033
rect -34 -347093 34 -347059
rect -34 -347201 34 -347167
rect -96 -348227 -62 -347251
rect 62 -348227 96 -347251
rect -34 -348311 34 -348277
rect -34 -348419 34 -348385
rect -96 -349445 -62 -348469
rect 62 -349445 96 -348469
rect -34 -349529 34 -349495
rect -34 -349637 34 -349603
rect -96 -350663 -62 -349687
rect 62 -350663 96 -349687
rect -34 -350747 34 -350713
rect -34 -350855 34 -350821
rect -96 -351881 -62 -350905
rect 62 -351881 96 -350905
rect -34 -351965 34 -351931
rect -34 -352073 34 -352039
rect -96 -353099 -62 -352123
rect 62 -353099 96 -352123
rect -34 -353183 34 -353149
rect -34 -353291 34 -353257
rect -96 -354317 -62 -353341
rect 62 -354317 96 -353341
rect -34 -354401 34 -354367
rect -34 -354509 34 -354475
rect -96 -355535 -62 -354559
rect 62 -355535 96 -354559
rect -34 -355619 34 -355585
rect -34 -355727 34 -355693
rect -96 -356753 -62 -355777
rect 62 -356753 96 -355777
rect -34 -356837 34 -356803
rect -34 -356945 34 -356911
rect -96 -357971 -62 -356995
rect 62 -357971 96 -356995
rect -34 -358055 34 -358021
rect -34 -358163 34 -358129
rect -96 -359189 -62 -358213
rect 62 -359189 96 -358213
rect -34 -359273 34 -359239
rect -34 -359381 34 -359347
rect -96 -360407 -62 -359431
rect 62 -360407 96 -359431
rect -34 -360491 34 -360457
rect -34 -360599 34 -360565
rect -96 -361625 -62 -360649
rect 62 -361625 96 -360649
rect -34 -361709 34 -361675
rect -34 -361817 34 -361783
rect -96 -362843 -62 -361867
rect 62 -362843 96 -361867
rect -34 -362927 34 -362893
rect -34 -363035 34 -363001
rect -96 -364061 -62 -363085
rect 62 -364061 96 -363085
rect -34 -364145 34 -364111
rect -34 -364253 34 -364219
rect -96 -365279 -62 -364303
rect 62 -365279 96 -364303
rect -34 -365363 34 -365329
rect -34 -365471 34 -365437
rect -96 -366497 -62 -365521
rect 62 -366497 96 -365521
rect -34 -366581 34 -366547
rect -34 -366689 34 -366655
rect -96 -367715 -62 -366739
rect 62 -367715 96 -366739
rect -34 -367799 34 -367765
rect -34 -367907 34 -367873
rect -96 -368933 -62 -367957
rect 62 -368933 96 -367957
rect -34 -369017 34 -368983
rect -34 -369125 34 -369091
rect -96 -370151 -62 -369175
rect 62 -370151 96 -369175
rect -34 -370235 34 -370201
rect -34 -370343 34 -370309
rect -96 -371369 -62 -370393
rect 62 -371369 96 -370393
rect -34 -371453 34 -371419
rect -34 -371561 34 -371527
rect -96 -372587 -62 -371611
rect 62 -372587 96 -371611
rect -34 -372671 34 -372637
rect -34 -372779 34 -372745
rect -96 -373805 -62 -372829
rect 62 -373805 96 -372829
rect -34 -373889 34 -373855
rect -34 -373997 34 -373963
rect -96 -375023 -62 -374047
rect 62 -375023 96 -374047
rect -34 -375107 34 -375073
rect -34 -375215 34 -375181
rect -96 -376241 -62 -375265
rect 62 -376241 96 -375265
rect -34 -376325 34 -376291
rect -34 -376433 34 -376399
rect -96 -377459 -62 -376483
rect 62 -377459 96 -376483
rect -34 -377543 34 -377509
rect -34 -377651 34 -377617
rect -96 -378677 -62 -377701
rect 62 -378677 96 -377701
rect -34 -378761 34 -378727
rect -34 -378869 34 -378835
rect -96 -379895 -62 -378919
rect 62 -379895 96 -378919
rect -34 -379979 34 -379945
rect -34 -380087 34 -380053
rect -96 -381113 -62 -380137
rect 62 -381113 96 -380137
rect -34 -381197 34 -381163
rect -34 -381305 34 -381271
rect -96 -382331 -62 -381355
rect 62 -382331 96 -381355
rect -34 -382415 34 -382381
rect -34 -382523 34 -382489
rect -96 -383549 -62 -382573
rect 62 -383549 96 -382573
rect -34 -383633 34 -383599
rect -34 -383741 34 -383707
rect -96 -384767 -62 -383791
rect 62 -384767 96 -383791
rect -34 -384851 34 -384817
rect -34 -384959 34 -384925
rect -96 -385985 -62 -385009
rect 62 -385985 96 -385009
rect -34 -386069 34 -386035
rect -34 -386177 34 -386143
rect -96 -387203 -62 -386227
rect 62 -387203 96 -386227
rect -34 -387287 34 -387253
rect -34 -387395 34 -387361
rect -96 -388421 -62 -387445
rect 62 -388421 96 -387445
rect -34 -388505 34 -388471
rect -34 -388613 34 -388579
rect -96 -389639 -62 -388663
rect 62 -389639 96 -388663
rect -34 -389723 34 -389689
rect -34 -389831 34 -389797
rect -96 -390857 -62 -389881
rect 62 -390857 96 -389881
rect -34 -390941 34 -390907
rect -34 -391049 34 -391015
rect -96 -392075 -62 -391099
rect 62 -392075 96 -391099
rect -34 -392159 34 -392125
rect -34 -392267 34 -392233
rect -96 -393293 -62 -392317
rect 62 -393293 96 -392317
rect -34 -393377 34 -393343
rect -34 -393485 34 -393451
rect -96 -394511 -62 -393535
rect 62 -394511 96 -393535
rect -34 -394595 34 -394561
rect -34 -394703 34 -394669
rect -96 -395729 -62 -394753
rect 62 -395729 96 -394753
rect -34 -395813 34 -395779
rect -34 -395921 34 -395887
rect -96 -396947 -62 -395971
rect 62 -396947 96 -395971
rect -34 -397031 34 -396997
rect -34 -397139 34 -397105
rect -96 -398165 -62 -397189
rect 62 -398165 96 -397189
rect -34 -398249 34 -398215
rect -34 -398357 34 -398323
rect -96 -399383 -62 -398407
rect 62 -399383 96 -398407
rect -34 -399467 34 -399433
rect -34 -399575 34 -399541
rect -96 -400601 -62 -399625
rect 62 -400601 96 -399625
rect -34 -400685 34 -400651
rect -34 -400793 34 -400759
rect -96 -401819 -62 -400843
rect 62 -401819 96 -400843
rect -34 -401903 34 -401869
rect -34 -402011 34 -401977
rect -96 -403037 -62 -402061
rect 62 -403037 96 -402061
rect -34 -403121 34 -403087
rect -34 -403229 34 -403195
rect -96 -404255 -62 -403279
rect 62 -404255 96 -403279
rect -34 -404339 34 -404305
rect -34 -404447 34 -404413
rect -96 -405473 -62 -404497
rect 62 -405473 96 -404497
rect -34 -405557 34 -405523
rect -34 -405665 34 -405631
rect -96 -406691 -62 -405715
rect 62 -406691 96 -405715
rect -34 -406775 34 -406741
rect -34 -406883 34 -406849
rect -96 -407909 -62 -406933
rect 62 -407909 96 -406933
rect -34 -407993 34 -407959
rect -34 -408101 34 -408067
rect -96 -409127 -62 -408151
rect 62 -409127 96 -408151
rect -34 -409211 34 -409177
rect -34 -409319 34 -409285
rect -96 -410345 -62 -409369
rect 62 -410345 96 -409369
rect -34 -410429 34 -410395
rect -34 -410537 34 -410503
rect -96 -411563 -62 -410587
rect 62 -411563 96 -410587
rect -34 -411647 34 -411613
rect -34 -411755 34 -411721
rect -96 -412781 -62 -411805
rect 62 -412781 96 -411805
rect -34 -412865 34 -412831
rect -34 -412973 34 -412939
rect -96 -413999 -62 -413023
rect 62 -413999 96 -413023
rect -34 -414083 34 -414049
rect -34 -414191 34 -414157
rect -96 -415217 -62 -414241
rect 62 -415217 96 -414241
rect -34 -415301 34 -415267
rect -34 -415409 34 -415375
rect -96 -416435 -62 -415459
rect 62 -416435 96 -415459
rect -34 -416519 34 -416485
rect -34 -416627 34 -416593
rect -96 -417653 -62 -416677
rect 62 -417653 96 -416677
rect -34 -417737 34 -417703
rect -34 -417845 34 -417811
rect -96 -418871 -62 -417895
rect 62 -418871 96 -417895
rect -34 -418955 34 -418921
rect -34 -419063 34 -419029
rect -96 -420089 -62 -419113
rect 62 -420089 96 -419113
rect -34 -420173 34 -420139
rect -34 -420281 34 -420247
rect -96 -421307 -62 -420331
rect 62 -421307 96 -420331
rect -34 -421391 34 -421357
rect -34 -421499 34 -421465
rect -96 -422525 -62 -421549
rect 62 -422525 96 -421549
rect -34 -422609 34 -422575
rect -34 -422717 34 -422683
rect -96 -423743 -62 -422767
rect 62 -423743 96 -422767
rect -34 -423827 34 -423793
rect -34 -423935 34 -423901
rect -96 -424961 -62 -423985
rect 62 -424961 96 -423985
rect -34 -425045 34 -425011
rect -34 -425153 34 -425119
rect -96 -426179 -62 -425203
rect 62 -426179 96 -425203
rect -34 -426263 34 -426229
rect -34 -426371 34 -426337
rect -96 -427397 -62 -426421
rect 62 -427397 96 -426421
rect -34 -427481 34 -427447
rect -34 -427589 34 -427555
rect -96 -428615 -62 -427639
rect 62 -428615 96 -427639
rect -34 -428699 34 -428665
rect -34 -428807 34 -428773
rect -96 -429833 -62 -428857
rect 62 -429833 96 -428857
rect -34 -429917 34 -429883
rect -34 -430025 34 -429991
rect -96 -431051 -62 -430075
rect 62 -431051 96 -430075
rect -34 -431135 34 -431101
rect -34 -431243 34 -431209
rect -96 -432269 -62 -431293
rect 62 -432269 96 -431293
rect -34 -432353 34 -432319
rect -34 -432461 34 -432427
rect -96 -433487 -62 -432511
rect 62 -433487 96 -432511
rect -34 -433571 34 -433537
rect -34 -433679 34 -433645
rect -96 -434705 -62 -433729
rect 62 -434705 96 -433729
rect -34 -434789 34 -434755
rect -34 -434897 34 -434863
rect -96 -435923 -62 -434947
rect 62 -435923 96 -434947
rect -34 -436007 34 -435973
rect -34 -436115 34 -436081
rect -96 -437141 -62 -436165
rect 62 -437141 96 -436165
rect -34 -437225 34 -437191
rect -34 -437333 34 -437299
rect -96 -438359 -62 -437383
rect 62 -438359 96 -437383
rect -34 -438443 34 -438409
rect -34 -438551 34 -438517
rect -96 -439577 -62 -438601
rect 62 -439577 96 -438601
rect -34 -439661 34 -439627
rect -34 -439769 34 -439735
rect -96 -440795 -62 -439819
rect 62 -440795 96 -439819
rect -34 -440879 34 -440845
rect -34 -440987 34 -440953
rect -96 -442013 -62 -441037
rect 62 -442013 96 -441037
rect -34 -442097 34 -442063
rect -34 -442205 34 -442171
rect -96 -443231 -62 -442255
rect 62 -443231 96 -442255
rect -34 -443315 34 -443281
rect -34 -443423 34 -443389
rect -96 -444449 -62 -443473
rect 62 -444449 96 -443473
rect -34 -444533 34 -444499
rect -34 -444641 34 -444607
rect -96 -445667 -62 -444691
rect 62 -445667 96 -444691
rect -34 -445751 34 -445717
rect -34 -445859 34 -445825
rect -96 -446885 -62 -445909
rect 62 -446885 96 -445909
rect -34 -446969 34 -446935
rect -34 -447077 34 -447043
rect -96 -448103 -62 -447127
rect 62 -448103 96 -447127
rect -34 -448187 34 -448153
rect -34 -448295 34 -448261
rect -96 -449321 -62 -448345
rect 62 -449321 96 -448345
rect -34 -449405 34 -449371
rect -34 -449513 34 -449479
rect -96 -450539 -62 -449563
rect 62 -450539 96 -449563
rect -34 -450623 34 -450589
rect -34 -450731 34 -450697
rect -96 -451757 -62 -450781
rect 62 -451757 96 -450781
rect -34 -451841 34 -451807
rect -34 -451949 34 -451915
rect -96 -452975 -62 -451999
rect 62 -452975 96 -451999
rect -34 -453059 34 -453025
rect -34 -453167 34 -453133
rect -96 -454193 -62 -453217
rect 62 -454193 96 -453217
rect -34 -454277 34 -454243
rect -34 -454385 34 -454351
rect -96 -455411 -62 -454435
rect 62 -455411 96 -454435
rect -34 -455495 34 -455461
rect -34 -455603 34 -455569
rect -96 -456629 -62 -455653
rect 62 -456629 96 -455653
rect -34 -456713 34 -456679
rect -34 -456821 34 -456787
rect -96 -457847 -62 -456871
rect 62 -457847 96 -456871
rect -34 -457931 34 -457897
rect -34 -458039 34 -458005
rect -96 -459065 -62 -458089
rect 62 -459065 96 -458089
rect -34 -459149 34 -459115
rect -34 -459257 34 -459223
rect -96 -460283 -62 -459307
rect 62 -460283 96 -459307
rect -34 -460367 34 -460333
rect -34 -460475 34 -460441
rect -96 -461501 -62 -460525
rect 62 -461501 96 -460525
rect -34 -461585 34 -461551
rect -34 -461693 34 -461659
rect -96 -462719 -62 -461743
rect 62 -462719 96 -461743
rect -34 -462803 34 -462769
rect -34 -462911 34 -462877
rect -96 -463937 -62 -462961
rect 62 -463937 96 -462961
rect -34 -464021 34 -463987
rect -34 -464129 34 -464095
rect -96 -465155 -62 -464179
rect 62 -465155 96 -464179
rect -34 -465239 34 -465205
rect -34 -465347 34 -465313
rect -96 -466373 -62 -465397
rect 62 -466373 96 -465397
rect -34 -466457 34 -466423
rect -34 -466565 34 -466531
rect -96 -467591 -62 -466615
rect 62 -467591 96 -466615
rect -34 -467675 34 -467641
rect -34 -467783 34 -467749
rect -96 -468809 -62 -467833
rect 62 -468809 96 -467833
rect -34 -468893 34 -468859
rect -34 -469001 34 -468967
rect -96 -470027 -62 -469051
rect 62 -470027 96 -469051
rect -34 -470111 34 -470077
rect -34 -470219 34 -470185
rect -96 -471245 -62 -470269
rect 62 -471245 96 -470269
rect -34 -471329 34 -471295
rect -34 -471437 34 -471403
rect -96 -472463 -62 -471487
rect 62 -472463 96 -471487
rect -34 -472547 34 -472513
rect -34 -472655 34 -472621
rect -96 -473681 -62 -472705
rect 62 -473681 96 -472705
rect -34 -473765 34 -473731
rect -34 -473873 34 -473839
rect -96 -474899 -62 -473923
rect 62 -474899 96 -473923
rect -34 -474983 34 -474949
rect -34 -475091 34 -475057
rect -96 -476117 -62 -475141
rect 62 -476117 96 -475141
rect -34 -476201 34 -476167
rect -34 -476309 34 -476275
rect -96 -477335 -62 -476359
rect 62 -477335 96 -476359
rect -34 -477419 34 -477385
rect -34 -477527 34 -477493
rect -96 -478553 -62 -477577
rect 62 -478553 96 -477577
rect -34 -478637 34 -478603
rect -34 -478745 34 -478711
rect -96 -479771 -62 -478795
rect 62 -479771 96 -478795
rect -34 -479855 34 -479821
rect -34 -479963 34 -479929
rect -96 -480989 -62 -480013
rect 62 -480989 96 -480013
rect -34 -481073 34 -481039
rect -34 -481181 34 -481147
rect -96 -482207 -62 -481231
rect 62 -482207 96 -481231
rect -34 -482291 34 -482257
rect -34 -482399 34 -482365
rect -96 -483425 -62 -482449
rect 62 -483425 96 -482449
rect -34 -483509 34 -483475
rect -34 -483617 34 -483583
rect -96 -484643 -62 -483667
rect 62 -484643 96 -483667
rect -34 -484727 34 -484693
rect -34 -484835 34 -484801
rect -96 -485861 -62 -484885
rect 62 -485861 96 -484885
rect -34 -485945 34 -485911
rect -34 -486053 34 -486019
rect -96 -487079 -62 -486103
rect 62 -487079 96 -486103
rect -34 -487163 34 -487129
rect -34 -487271 34 -487237
rect -96 -488297 -62 -487321
rect 62 -488297 96 -487321
rect -34 -488381 34 -488347
rect -34 -488489 34 -488455
rect -96 -489515 -62 -488539
rect 62 -489515 96 -488539
rect -34 -489599 34 -489565
rect -34 -489707 34 -489673
rect -96 -490733 -62 -489757
rect 62 -490733 96 -489757
rect -34 -490817 34 -490783
rect -34 -490925 34 -490891
rect -96 -491951 -62 -490975
rect 62 -491951 96 -490975
rect -34 -492035 34 -492001
rect -34 -492143 34 -492109
rect -96 -493169 -62 -492193
rect 62 -493169 96 -492193
rect -34 -493253 34 -493219
rect -34 -493361 34 -493327
rect -96 -494387 -62 -493411
rect 62 -494387 96 -493411
rect -34 -494471 34 -494437
rect -34 -494579 34 -494545
rect -96 -495605 -62 -494629
rect 62 -495605 96 -494629
rect -34 -495689 34 -495655
rect -34 -495797 34 -495763
rect -96 -496823 -62 -495847
rect 62 -496823 96 -495847
rect -34 -496907 34 -496873
rect -34 -497015 34 -496981
rect -96 -498041 -62 -497065
rect 62 -498041 96 -497065
rect -34 -498125 34 -498091
rect -34 -498233 34 -498199
rect -96 -499259 -62 -498283
rect 62 -499259 96 -498283
rect -34 -499343 34 -499309
rect -34 -499451 34 -499417
rect -96 -500477 -62 -499501
rect 62 -500477 96 -499501
rect -34 -500561 34 -500527
rect -34 -500669 34 -500635
rect -96 -501695 -62 -500719
rect 62 -501695 96 -500719
rect -34 -501779 34 -501745
rect -34 -501887 34 -501853
rect -96 -502913 -62 -501937
rect 62 -502913 96 -501937
rect -34 -502997 34 -502963
rect -34 -503105 34 -503071
rect -96 -504131 -62 -503155
rect 62 -504131 96 -503155
rect -34 -504215 34 -504181
rect -34 -504323 34 -504289
rect -96 -505349 -62 -504373
rect 62 -505349 96 -504373
rect -34 -505433 34 -505399
rect -34 -505541 34 -505507
rect -96 -506567 -62 -505591
rect 62 -506567 96 -505591
rect -34 -506651 34 -506617
rect -34 -506759 34 -506725
rect -96 -507785 -62 -506809
rect 62 -507785 96 -506809
rect -34 -507869 34 -507835
rect -34 -507977 34 -507943
rect -96 -509003 -62 -508027
rect 62 -509003 96 -508027
rect -34 -509087 34 -509053
rect -34 -509195 34 -509161
rect -96 -510221 -62 -509245
rect 62 -510221 96 -509245
rect -34 -510305 34 -510271
rect -34 -510413 34 -510379
rect -96 -511439 -62 -510463
rect 62 -511439 96 -510463
rect -34 -511523 34 -511489
rect -34 -511631 34 -511597
rect -96 -512657 -62 -511681
rect 62 -512657 96 -511681
rect -34 -512741 34 -512707
rect -34 -512849 34 -512815
rect -96 -513875 -62 -512899
rect 62 -513875 96 -512899
rect -34 -513959 34 -513925
rect -34 -514067 34 -514033
rect -96 -515093 -62 -514117
rect 62 -515093 96 -514117
rect -34 -515177 34 -515143
rect -34 -515285 34 -515251
rect -96 -516311 -62 -515335
rect 62 -516311 96 -515335
rect -34 -516395 34 -516361
rect -34 -516503 34 -516469
rect -96 -517529 -62 -516553
rect 62 -517529 96 -516553
rect -34 -517613 34 -517579
rect -34 -517721 34 -517687
rect -96 -518747 -62 -517771
rect 62 -518747 96 -517771
rect -34 -518831 34 -518797
rect -34 -518939 34 -518905
rect -96 -519965 -62 -518989
rect 62 -519965 96 -518989
rect -34 -520049 34 -520015
rect -34 -520157 34 -520123
rect -96 -521183 -62 -520207
rect 62 -521183 96 -520207
rect -34 -521267 34 -521233
rect -34 -521375 34 -521341
rect -96 -522401 -62 -521425
rect 62 -522401 96 -521425
rect -34 -522485 34 -522451
rect -34 -522593 34 -522559
rect -96 -523619 -62 -522643
rect 62 -523619 96 -522643
rect -34 -523703 34 -523669
rect -34 -523811 34 -523777
rect -96 -524837 -62 -523861
rect 62 -524837 96 -523861
rect -34 -524921 34 -524887
rect -34 -525029 34 -524995
rect -96 -526055 -62 -525079
rect 62 -526055 96 -525079
rect -34 -526139 34 -526105
rect -34 -526247 34 -526213
rect -96 -527273 -62 -526297
rect 62 -527273 96 -526297
rect -34 -527357 34 -527323
rect -34 -527465 34 -527431
rect -96 -528491 -62 -527515
rect 62 -528491 96 -527515
rect -34 -528575 34 -528541
rect -34 -528683 34 -528649
rect -96 -529709 -62 -528733
rect 62 -529709 96 -528733
rect -34 -529793 34 -529759
rect -34 -529901 34 -529867
rect -96 -530927 -62 -529951
rect 62 -530927 96 -529951
rect -34 -531011 34 -530977
rect -34 -531119 34 -531085
rect -96 -532145 -62 -531169
rect 62 -532145 96 -531169
rect -34 -532229 34 -532195
rect -34 -532337 34 -532303
rect -96 -533363 -62 -532387
rect 62 -533363 96 -532387
rect -34 -533447 34 -533413
rect -34 -533555 34 -533521
rect -96 -534581 -62 -533605
rect 62 -534581 96 -533605
rect -34 -534665 34 -534631
rect -34 -534773 34 -534739
rect -96 -535799 -62 -534823
rect 62 -535799 96 -534823
rect -34 -535883 34 -535849
rect -34 -535991 34 -535957
rect -96 -537017 -62 -536041
rect 62 -537017 96 -536041
rect -34 -537101 34 -537067
rect -34 -537209 34 -537175
rect -96 -538235 -62 -537259
rect 62 -538235 96 -537259
rect -34 -538319 34 -538285
rect -34 -538427 34 -538393
rect -96 -539453 -62 -538477
rect 62 -539453 96 -538477
rect -34 -539537 34 -539503
rect -34 -539645 34 -539611
rect -96 -540671 -62 -539695
rect 62 -540671 96 -539695
rect -34 -540755 34 -540721
rect -34 -540863 34 -540829
rect -96 -541889 -62 -540913
rect 62 -541889 96 -540913
rect -34 -541973 34 -541939
rect -34 -542081 34 -542047
rect -96 -543107 -62 -542131
rect 62 -543107 96 -542131
rect -34 -543191 34 -543157
rect -34 -543299 34 -543265
rect -96 -544325 -62 -543349
rect 62 -544325 96 -543349
rect -34 -544409 34 -544375
rect -34 -544517 34 -544483
rect -96 -545543 -62 -544567
rect 62 -545543 96 -544567
rect -34 -545627 34 -545593
rect -34 -545735 34 -545701
rect -96 -546761 -62 -545785
rect 62 -546761 96 -545785
rect -34 -546845 34 -546811
rect -34 -546953 34 -546919
rect -96 -547979 -62 -547003
rect 62 -547979 96 -547003
rect -34 -548063 34 -548029
rect -34 -548171 34 -548137
rect -96 -549197 -62 -548221
rect 62 -549197 96 -548221
rect -34 -549281 34 -549247
rect -34 -549389 34 -549355
rect -96 -550415 -62 -549439
rect 62 -550415 96 -549439
rect -34 -550499 34 -550465
rect -34 -550607 34 -550573
rect -96 -551633 -62 -550657
rect 62 -551633 96 -550657
rect -34 -551717 34 -551683
rect -34 -551825 34 -551791
rect -96 -552851 -62 -551875
rect 62 -552851 96 -551875
rect -34 -552935 34 -552901
rect -34 -553043 34 -553009
rect -96 -554069 -62 -553093
rect 62 -554069 96 -553093
rect -34 -554153 34 -554119
rect -34 -554261 34 -554227
rect -96 -555287 -62 -554311
rect 62 -555287 96 -554311
rect -34 -555371 34 -555337
rect -34 -555479 34 -555445
rect -96 -556505 -62 -555529
rect 62 -556505 96 -555529
rect -34 -556589 34 -556555
rect -34 -556697 34 -556663
rect -96 -557723 -62 -556747
rect 62 -557723 96 -556747
rect -34 -557807 34 -557773
rect -34 -557915 34 -557881
rect -96 -558941 -62 -557965
rect 62 -558941 96 -557965
rect -34 -559025 34 -558991
rect -34 -559133 34 -559099
rect -96 -560159 -62 -559183
rect 62 -560159 96 -559183
rect -34 -560243 34 -560209
rect -34 -560351 34 -560317
rect -96 -561377 -62 -560401
rect 62 -561377 96 -560401
rect -34 -561461 34 -561427
rect -34 -561569 34 -561535
rect -96 -562595 -62 -561619
rect 62 -562595 96 -561619
rect -34 -562679 34 -562645
rect -34 -562787 34 -562753
rect -96 -563813 -62 -562837
rect 62 -563813 96 -562837
rect -34 -563897 34 -563863
rect -34 -564005 34 -563971
rect -96 -565031 -62 -564055
rect 62 -565031 96 -564055
rect -34 -565115 34 -565081
rect -34 -565223 34 -565189
rect -96 -566249 -62 -565273
rect 62 -566249 96 -565273
rect -34 -566333 34 -566299
rect -34 -566441 34 -566407
rect -96 -567467 -62 -566491
rect 62 -567467 96 -566491
rect -34 -567551 34 -567517
rect -34 -567659 34 -567625
rect -96 -568685 -62 -567709
rect 62 -568685 96 -567709
rect -34 -568769 34 -568735
rect -34 -568877 34 -568843
rect -96 -569903 -62 -568927
rect 62 -569903 96 -568927
rect -34 -569987 34 -569953
rect -34 -570095 34 -570061
rect -96 -571121 -62 -570145
rect 62 -571121 96 -570145
rect -34 -571205 34 -571171
rect -34 -571313 34 -571279
rect -96 -572339 -62 -571363
rect 62 -572339 96 -571363
rect -34 -572423 34 -572389
rect -34 -572531 34 -572497
rect -96 -573557 -62 -572581
rect 62 -573557 96 -572581
rect -34 -573641 34 -573607
rect -34 -573749 34 -573715
rect -96 -574775 -62 -573799
rect 62 -574775 96 -573799
rect -34 -574859 34 -574825
rect -34 -574967 34 -574933
rect -96 -575993 -62 -575017
rect 62 -575993 96 -575017
rect -34 -576077 34 -576043
rect -34 -576185 34 -576151
rect -96 -577211 -62 -576235
rect 62 -577211 96 -576235
rect -34 -577295 34 -577261
rect -34 -577403 34 -577369
rect -96 -578429 -62 -577453
rect 62 -578429 96 -577453
rect -34 -578513 34 -578479
rect -34 -578621 34 -578587
rect -96 -579647 -62 -578671
rect 62 -579647 96 -578671
rect -34 -579731 34 -579697
rect -34 -579839 34 -579805
rect -96 -580865 -62 -579889
rect 62 -580865 96 -579889
rect -34 -580949 34 -580915
rect -34 -581057 34 -581023
rect -96 -582083 -62 -581107
rect 62 -582083 96 -581107
rect -34 -582167 34 -582133
rect -34 -582275 34 -582241
rect -96 -583301 -62 -582325
rect 62 -583301 96 -582325
rect -34 -583385 34 -583351
rect -34 -583493 34 -583459
rect -96 -584519 -62 -583543
rect 62 -584519 96 -583543
rect -34 -584603 34 -584569
rect -34 -584711 34 -584677
rect -96 -585737 -62 -584761
rect 62 -585737 96 -584761
rect -34 -585821 34 -585787
rect -34 -585929 34 -585895
rect -96 -586955 -62 -585979
rect 62 -586955 96 -585979
rect -34 -587039 34 -587005
rect -34 -587147 34 -587113
rect -96 -588173 -62 -587197
rect 62 -588173 96 -587197
rect -34 -588257 34 -588223
rect -34 -588365 34 -588331
rect -96 -589391 -62 -588415
rect 62 -589391 96 -588415
rect -34 -589475 34 -589441
rect -34 -589583 34 -589549
rect -96 -590609 -62 -589633
rect 62 -590609 96 -589633
rect -34 -590693 34 -590659
rect -34 -590801 34 -590767
rect -96 -591827 -62 -590851
rect 62 -591827 96 -590851
rect -34 -591911 34 -591877
rect -34 -592019 34 -591985
rect -96 -593045 -62 -592069
rect 62 -593045 96 -592069
rect -34 -593129 34 -593095
rect -34 -593237 34 -593203
rect -96 -594263 -62 -593287
rect 62 -594263 96 -593287
rect -34 -594347 34 -594313
rect -34 -594455 34 -594421
rect -96 -595481 -62 -594505
rect 62 -595481 96 -594505
rect -34 -595565 34 -595531
rect -34 -595673 34 -595639
rect -96 -596699 -62 -595723
rect 62 -596699 96 -595723
rect -34 -596783 34 -596749
rect -34 -596891 34 -596857
rect -96 -597917 -62 -596941
rect 62 -597917 96 -596941
rect -34 -598001 34 -597967
rect -34 -598109 34 -598075
rect -96 -599135 -62 -598159
rect 62 -599135 96 -598159
rect -34 -599219 34 -599185
rect -34 -599327 34 -599293
rect -96 -600353 -62 -599377
rect 62 -600353 96 -599377
rect -34 -600437 34 -600403
rect -34 -600545 34 -600511
rect -96 -601571 -62 -600595
rect 62 -601571 96 -600595
rect -34 -601655 34 -601621
rect -34 -601763 34 -601729
rect -96 -602789 -62 -601813
rect 62 -602789 96 -601813
rect -34 -602873 34 -602839
rect -34 -602981 34 -602947
rect -96 -604007 -62 -603031
rect 62 -604007 96 -603031
rect -34 -604091 34 -604057
rect -34 -604199 34 -604165
rect -96 -605225 -62 -604249
rect 62 -605225 96 -604249
rect -34 -605309 34 -605275
rect -34 -605417 34 -605383
rect -96 -606443 -62 -605467
rect 62 -606443 96 -605467
rect -34 -606527 34 -606493
rect -34 -606635 34 -606601
rect -96 -607661 -62 -606685
rect 62 -607661 96 -606685
rect -34 -607745 34 -607711
rect -34 -607853 34 -607819
rect -96 -608879 -62 -607903
rect 62 -608879 96 -607903
rect -34 -608963 34 -608929
<< metal1 >>
rect -46 608963 46 608969
rect -46 608929 -34 608963
rect 34 608929 46 608963
rect -46 608923 46 608929
rect -102 608879 -56 608891
rect -102 607903 -96 608879
rect -62 607903 -56 608879
rect -102 607891 -56 607903
rect 56 608879 102 608891
rect 56 607903 62 608879
rect 96 607903 102 608879
rect 56 607891 102 607903
rect -46 607853 46 607859
rect -46 607819 -34 607853
rect 34 607819 46 607853
rect -46 607813 46 607819
rect -46 607745 46 607751
rect -46 607711 -34 607745
rect 34 607711 46 607745
rect -46 607705 46 607711
rect -102 607661 -56 607673
rect -102 606685 -96 607661
rect -62 606685 -56 607661
rect -102 606673 -56 606685
rect 56 607661 102 607673
rect 56 606685 62 607661
rect 96 606685 102 607661
rect 56 606673 102 606685
rect -46 606635 46 606641
rect -46 606601 -34 606635
rect 34 606601 46 606635
rect -46 606595 46 606601
rect -46 606527 46 606533
rect -46 606493 -34 606527
rect 34 606493 46 606527
rect -46 606487 46 606493
rect -102 606443 -56 606455
rect -102 605467 -96 606443
rect -62 605467 -56 606443
rect -102 605455 -56 605467
rect 56 606443 102 606455
rect 56 605467 62 606443
rect 96 605467 102 606443
rect 56 605455 102 605467
rect -46 605417 46 605423
rect -46 605383 -34 605417
rect 34 605383 46 605417
rect -46 605377 46 605383
rect -46 605309 46 605315
rect -46 605275 -34 605309
rect 34 605275 46 605309
rect -46 605269 46 605275
rect -102 605225 -56 605237
rect -102 604249 -96 605225
rect -62 604249 -56 605225
rect -102 604237 -56 604249
rect 56 605225 102 605237
rect 56 604249 62 605225
rect 96 604249 102 605225
rect 56 604237 102 604249
rect -46 604199 46 604205
rect -46 604165 -34 604199
rect 34 604165 46 604199
rect -46 604159 46 604165
rect -46 604091 46 604097
rect -46 604057 -34 604091
rect 34 604057 46 604091
rect -46 604051 46 604057
rect -102 604007 -56 604019
rect -102 603031 -96 604007
rect -62 603031 -56 604007
rect -102 603019 -56 603031
rect 56 604007 102 604019
rect 56 603031 62 604007
rect 96 603031 102 604007
rect 56 603019 102 603031
rect -46 602981 46 602987
rect -46 602947 -34 602981
rect 34 602947 46 602981
rect -46 602941 46 602947
rect -46 602873 46 602879
rect -46 602839 -34 602873
rect 34 602839 46 602873
rect -46 602833 46 602839
rect -102 602789 -56 602801
rect -102 601813 -96 602789
rect -62 601813 -56 602789
rect -102 601801 -56 601813
rect 56 602789 102 602801
rect 56 601813 62 602789
rect 96 601813 102 602789
rect 56 601801 102 601813
rect -46 601763 46 601769
rect -46 601729 -34 601763
rect 34 601729 46 601763
rect -46 601723 46 601729
rect -46 601655 46 601661
rect -46 601621 -34 601655
rect 34 601621 46 601655
rect -46 601615 46 601621
rect -102 601571 -56 601583
rect -102 600595 -96 601571
rect -62 600595 -56 601571
rect -102 600583 -56 600595
rect 56 601571 102 601583
rect 56 600595 62 601571
rect 96 600595 102 601571
rect 56 600583 102 600595
rect -46 600545 46 600551
rect -46 600511 -34 600545
rect 34 600511 46 600545
rect -46 600505 46 600511
rect -46 600437 46 600443
rect -46 600403 -34 600437
rect 34 600403 46 600437
rect -46 600397 46 600403
rect -102 600353 -56 600365
rect -102 599377 -96 600353
rect -62 599377 -56 600353
rect -102 599365 -56 599377
rect 56 600353 102 600365
rect 56 599377 62 600353
rect 96 599377 102 600353
rect 56 599365 102 599377
rect -46 599327 46 599333
rect -46 599293 -34 599327
rect 34 599293 46 599327
rect -46 599287 46 599293
rect -46 599219 46 599225
rect -46 599185 -34 599219
rect 34 599185 46 599219
rect -46 599179 46 599185
rect -102 599135 -56 599147
rect -102 598159 -96 599135
rect -62 598159 -56 599135
rect -102 598147 -56 598159
rect 56 599135 102 599147
rect 56 598159 62 599135
rect 96 598159 102 599135
rect 56 598147 102 598159
rect -46 598109 46 598115
rect -46 598075 -34 598109
rect 34 598075 46 598109
rect -46 598069 46 598075
rect -46 598001 46 598007
rect -46 597967 -34 598001
rect 34 597967 46 598001
rect -46 597961 46 597967
rect -102 597917 -56 597929
rect -102 596941 -96 597917
rect -62 596941 -56 597917
rect -102 596929 -56 596941
rect 56 597917 102 597929
rect 56 596941 62 597917
rect 96 596941 102 597917
rect 56 596929 102 596941
rect -46 596891 46 596897
rect -46 596857 -34 596891
rect 34 596857 46 596891
rect -46 596851 46 596857
rect -46 596783 46 596789
rect -46 596749 -34 596783
rect 34 596749 46 596783
rect -46 596743 46 596749
rect -102 596699 -56 596711
rect -102 595723 -96 596699
rect -62 595723 -56 596699
rect -102 595711 -56 595723
rect 56 596699 102 596711
rect 56 595723 62 596699
rect 96 595723 102 596699
rect 56 595711 102 595723
rect -46 595673 46 595679
rect -46 595639 -34 595673
rect 34 595639 46 595673
rect -46 595633 46 595639
rect -46 595565 46 595571
rect -46 595531 -34 595565
rect 34 595531 46 595565
rect -46 595525 46 595531
rect -102 595481 -56 595493
rect -102 594505 -96 595481
rect -62 594505 -56 595481
rect -102 594493 -56 594505
rect 56 595481 102 595493
rect 56 594505 62 595481
rect 96 594505 102 595481
rect 56 594493 102 594505
rect -46 594455 46 594461
rect -46 594421 -34 594455
rect 34 594421 46 594455
rect -46 594415 46 594421
rect -46 594347 46 594353
rect -46 594313 -34 594347
rect 34 594313 46 594347
rect -46 594307 46 594313
rect -102 594263 -56 594275
rect -102 593287 -96 594263
rect -62 593287 -56 594263
rect -102 593275 -56 593287
rect 56 594263 102 594275
rect 56 593287 62 594263
rect 96 593287 102 594263
rect 56 593275 102 593287
rect -46 593237 46 593243
rect -46 593203 -34 593237
rect 34 593203 46 593237
rect -46 593197 46 593203
rect -46 593129 46 593135
rect -46 593095 -34 593129
rect 34 593095 46 593129
rect -46 593089 46 593095
rect -102 593045 -56 593057
rect -102 592069 -96 593045
rect -62 592069 -56 593045
rect -102 592057 -56 592069
rect 56 593045 102 593057
rect 56 592069 62 593045
rect 96 592069 102 593045
rect 56 592057 102 592069
rect -46 592019 46 592025
rect -46 591985 -34 592019
rect 34 591985 46 592019
rect -46 591979 46 591985
rect -46 591911 46 591917
rect -46 591877 -34 591911
rect 34 591877 46 591911
rect -46 591871 46 591877
rect -102 591827 -56 591839
rect -102 590851 -96 591827
rect -62 590851 -56 591827
rect -102 590839 -56 590851
rect 56 591827 102 591839
rect 56 590851 62 591827
rect 96 590851 102 591827
rect 56 590839 102 590851
rect -46 590801 46 590807
rect -46 590767 -34 590801
rect 34 590767 46 590801
rect -46 590761 46 590767
rect -46 590693 46 590699
rect -46 590659 -34 590693
rect 34 590659 46 590693
rect -46 590653 46 590659
rect -102 590609 -56 590621
rect -102 589633 -96 590609
rect -62 589633 -56 590609
rect -102 589621 -56 589633
rect 56 590609 102 590621
rect 56 589633 62 590609
rect 96 589633 102 590609
rect 56 589621 102 589633
rect -46 589583 46 589589
rect -46 589549 -34 589583
rect 34 589549 46 589583
rect -46 589543 46 589549
rect -46 589475 46 589481
rect -46 589441 -34 589475
rect 34 589441 46 589475
rect -46 589435 46 589441
rect -102 589391 -56 589403
rect -102 588415 -96 589391
rect -62 588415 -56 589391
rect -102 588403 -56 588415
rect 56 589391 102 589403
rect 56 588415 62 589391
rect 96 588415 102 589391
rect 56 588403 102 588415
rect -46 588365 46 588371
rect -46 588331 -34 588365
rect 34 588331 46 588365
rect -46 588325 46 588331
rect -46 588257 46 588263
rect -46 588223 -34 588257
rect 34 588223 46 588257
rect -46 588217 46 588223
rect -102 588173 -56 588185
rect -102 587197 -96 588173
rect -62 587197 -56 588173
rect -102 587185 -56 587197
rect 56 588173 102 588185
rect 56 587197 62 588173
rect 96 587197 102 588173
rect 56 587185 102 587197
rect -46 587147 46 587153
rect -46 587113 -34 587147
rect 34 587113 46 587147
rect -46 587107 46 587113
rect -46 587039 46 587045
rect -46 587005 -34 587039
rect 34 587005 46 587039
rect -46 586999 46 587005
rect -102 586955 -56 586967
rect -102 585979 -96 586955
rect -62 585979 -56 586955
rect -102 585967 -56 585979
rect 56 586955 102 586967
rect 56 585979 62 586955
rect 96 585979 102 586955
rect 56 585967 102 585979
rect -46 585929 46 585935
rect -46 585895 -34 585929
rect 34 585895 46 585929
rect -46 585889 46 585895
rect -46 585821 46 585827
rect -46 585787 -34 585821
rect 34 585787 46 585821
rect -46 585781 46 585787
rect -102 585737 -56 585749
rect -102 584761 -96 585737
rect -62 584761 -56 585737
rect -102 584749 -56 584761
rect 56 585737 102 585749
rect 56 584761 62 585737
rect 96 584761 102 585737
rect 56 584749 102 584761
rect -46 584711 46 584717
rect -46 584677 -34 584711
rect 34 584677 46 584711
rect -46 584671 46 584677
rect -46 584603 46 584609
rect -46 584569 -34 584603
rect 34 584569 46 584603
rect -46 584563 46 584569
rect -102 584519 -56 584531
rect -102 583543 -96 584519
rect -62 583543 -56 584519
rect -102 583531 -56 583543
rect 56 584519 102 584531
rect 56 583543 62 584519
rect 96 583543 102 584519
rect 56 583531 102 583543
rect -46 583493 46 583499
rect -46 583459 -34 583493
rect 34 583459 46 583493
rect -46 583453 46 583459
rect -46 583385 46 583391
rect -46 583351 -34 583385
rect 34 583351 46 583385
rect -46 583345 46 583351
rect -102 583301 -56 583313
rect -102 582325 -96 583301
rect -62 582325 -56 583301
rect -102 582313 -56 582325
rect 56 583301 102 583313
rect 56 582325 62 583301
rect 96 582325 102 583301
rect 56 582313 102 582325
rect -46 582275 46 582281
rect -46 582241 -34 582275
rect 34 582241 46 582275
rect -46 582235 46 582241
rect -46 582167 46 582173
rect -46 582133 -34 582167
rect 34 582133 46 582167
rect -46 582127 46 582133
rect -102 582083 -56 582095
rect -102 581107 -96 582083
rect -62 581107 -56 582083
rect -102 581095 -56 581107
rect 56 582083 102 582095
rect 56 581107 62 582083
rect 96 581107 102 582083
rect 56 581095 102 581107
rect -46 581057 46 581063
rect -46 581023 -34 581057
rect 34 581023 46 581057
rect -46 581017 46 581023
rect -46 580949 46 580955
rect -46 580915 -34 580949
rect 34 580915 46 580949
rect -46 580909 46 580915
rect -102 580865 -56 580877
rect -102 579889 -96 580865
rect -62 579889 -56 580865
rect -102 579877 -56 579889
rect 56 580865 102 580877
rect 56 579889 62 580865
rect 96 579889 102 580865
rect 56 579877 102 579889
rect -46 579839 46 579845
rect -46 579805 -34 579839
rect 34 579805 46 579839
rect -46 579799 46 579805
rect -46 579731 46 579737
rect -46 579697 -34 579731
rect 34 579697 46 579731
rect -46 579691 46 579697
rect -102 579647 -56 579659
rect -102 578671 -96 579647
rect -62 578671 -56 579647
rect -102 578659 -56 578671
rect 56 579647 102 579659
rect 56 578671 62 579647
rect 96 578671 102 579647
rect 56 578659 102 578671
rect -46 578621 46 578627
rect -46 578587 -34 578621
rect 34 578587 46 578621
rect -46 578581 46 578587
rect -46 578513 46 578519
rect -46 578479 -34 578513
rect 34 578479 46 578513
rect -46 578473 46 578479
rect -102 578429 -56 578441
rect -102 577453 -96 578429
rect -62 577453 -56 578429
rect -102 577441 -56 577453
rect 56 578429 102 578441
rect 56 577453 62 578429
rect 96 577453 102 578429
rect 56 577441 102 577453
rect -46 577403 46 577409
rect -46 577369 -34 577403
rect 34 577369 46 577403
rect -46 577363 46 577369
rect -46 577295 46 577301
rect -46 577261 -34 577295
rect 34 577261 46 577295
rect -46 577255 46 577261
rect -102 577211 -56 577223
rect -102 576235 -96 577211
rect -62 576235 -56 577211
rect -102 576223 -56 576235
rect 56 577211 102 577223
rect 56 576235 62 577211
rect 96 576235 102 577211
rect 56 576223 102 576235
rect -46 576185 46 576191
rect -46 576151 -34 576185
rect 34 576151 46 576185
rect -46 576145 46 576151
rect -46 576077 46 576083
rect -46 576043 -34 576077
rect 34 576043 46 576077
rect -46 576037 46 576043
rect -102 575993 -56 576005
rect -102 575017 -96 575993
rect -62 575017 -56 575993
rect -102 575005 -56 575017
rect 56 575993 102 576005
rect 56 575017 62 575993
rect 96 575017 102 575993
rect 56 575005 102 575017
rect -46 574967 46 574973
rect -46 574933 -34 574967
rect 34 574933 46 574967
rect -46 574927 46 574933
rect -46 574859 46 574865
rect -46 574825 -34 574859
rect 34 574825 46 574859
rect -46 574819 46 574825
rect -102 574775 -56 574787
rect -102 573799 -96 574775
rect -62 573799 -56 574775
rect -102 573787 -56 573799
rect 56 574775 102 574787
rect 56 573799 62 574775
rect 96 573799 102 574775
rect 56 573787 102 573799
rect -46 573749 46 573755
rect -46 573715 -34 573749
rect 34 573715 46 573749
rect -46 573709 46 573715
rect -46 573641 46 573647
rect -46 573607 -34 573641
rect 34 573607 46 573641
rect -46 573601 46 573607
rect -102 573557 -56 573569
rect -102 572581 -96 573557
rect -62 572581 -56 573557
rect -102 572569 -56 572581
rect 56 573557 102 573569
rect 56 572581 62 573557
rect 96 572581 102 573557
rect 56 572569 102 572581
rect -46 572531 46 572537
rect -46 572497 -34 572531
rect 34 572497 46 572531
rect -46 572491 46 572497
rect -46 572423 46 572429
rect -46 572389 -34 572423
rect 34 572389 46 572423
rect -46 572383 46 572389
rect -102 572339 -56 572351
rect -102 571363 -96 572339
rect -62 571363 -56 572339
rect -102 571351 -56 571363
rect 56 572339 102 572351
rect 56 571363 62 572339
rect 96 571363 102 572339
rect 56 571351 102 571363
rect -46 571313 46 571319
rect -46 571279 -34 571313
rect 34 571279 46 571313
rect -46 571273 46 571279
rect -46 571205 46 571211
rect -46 571171 -34 571205
rect 34 571171 46 571205
rect -46 571165 46 571171
rect -102 571121 -56 571133
rect -102 570145 -96 571121
rect -62 570145 -56 571121
rect -102 570133 -56 570145
rect 56 571121 102 571133
rect 56 570145 62 571121
rect 96 570145 102 571121
rect 56 570133 102 570145
rect -46 570095 46 570101
rect -46 570061 -34 570095
rect 34 570061 46 570095
rect -46 570055 46 570061
rect -46 569987 46 569993
rect -46 569953 -34 569987
rect 34 569953 46 569987
rect -46 569947 46 569953
rect -102 569903 -56 569915
rect -102 568927 -96 569903
rect -62 568927 -56 569903
rect -102 568915 -56 568927
rect 56 569903 102 569915
rect 56 568927 62 569903
rect 96 568927 102 569903
rect 56 568915 102 568927
rect -46 568877 46 568883
rect -46 568843 -34 568877
rect 34 568843 46 568877
rect -46 568837 46 568843
rect -46 568769 46 568775
rect -46 568735 -34 568769
rect 34 568735 46 568769
rect -46 568729 46 568735
rect -102 568685 -56 568697
rect -102 567709 -96 568685
rect -62 567709 -56 568685
rect -102 567697 -56 567709
rect 56 568685 102 568697
rect 56 567709 62 568685
rect 96 567709 102 568685
rect 56 567697 102 567709
rect -46 567659 46 567665
rect -46 567625 -34 567659
rect 34 567625 46 567659
rect -46 567619 46 567625
rect -46 567551 46 567557
rect -46 567517 -34 567551
rect 34 567517 46 567551
rect -46 567511 46 567517
rect -102 567467 -56 567479
rect -102 566491 -96 567467
rect -62 566491 -56 567467
rect -102 566479 -56 566491
rect 56 567467 102 567479
rect 56 566491 62 567467
rect 96 566491 102 567467
rect 56 566479 102 566491
rect -46 566441 46 566447
rect -46 566407 -34 566441
rect 34 566407 46 566441
rect -46 566401 46 566407
rect -46 566333 46 566339
rect -46 566299 -34 566333
rect 34 566299 46 566333
rect -46 566293 46 566299
rect -102 566249 -56 566261
rect -102 565273 -96 566249
rect -62 565273 -56 566249
rect -102 565261 -56 565273
rect 56 566249 102 566261
rect 56 565273 62 566249
rect 96 565273 102 566249
rect 56 565261 102 565273
rect -46 565223 46 565229
rect -46 565189 -34 565223
rect 34 565189 46 565223
rect -46 565183 46 565189
rect -46 565115 46 565121
rect -46 565081 -34 565115
rect 34 565081 46 565115
rect -46 565075 46 565081
rect -102 565031 -56 565043
rect -102 564055 -96 565031
rect -62 564055 -56 565031
rect -102 564043 -56 564055
rect 56 565031 102 565043
rect 56 564055 62 565031
rect 96 564055 102 565031
rect 56 564043 102 564055
rect -46 564005 46 564011
rect -46 563971 -34 564005
rect 34 563971 46 564005
rect -46 563965 46 563971
rect -46 563897 46 563903
rect -46 563863 -34 563897
rect 34 563863 46 563897
rect -46 563857 46 563863
rect -102 563813 -56 563825
rect -102 562837 -96 563813
rect -62 562837 -56 563813
rect -102 562825 -56 562837
rect 56 563813 102 563825
rect 56 562837 62 563813
rect 96 562837 102 563813
rect 56 562825 102 562837
rect -46 562787 46 562793
rect -46 562753 -34 562787
rect 34 562753 46 562787
rect -46 562747 46 562753
rect -46 562679 46 562685
rect -46 562645 -34 562679
rect 34 562645 46 562679
rect -46 562639 46 562645
rect -102 562595 -56 562607
rect -102 561619 -96 562595
rect -62 561619 -56 562595
rect -102 561607 -56 561619
rect 56 562595 102 562607
rect 56 561619 62 562595
rect 96 561619 102 562595
rect 56 561607 102 561619
rect -46 561569 46 561575
rect -46 561535 -34 561569
rect 34 561535 46 561569
rect -46 561529 46 561535
rect -46 561461 46 561467
rect -46 561427 -34 561461
rect 34 561427 46 561461
rect -46 561421 46 561427
rect -102 561377 -56 561389
rect -102 560401 -96 561377
rect -62 560401 -56 561377
rect -102 560389 -56 560401
rect 56 561377 102 561389
rect 56 560401 62 561377
rect 96 560401 102 561377
rect 56 560389 102 560401
rect -46 560351 46 560357
rect -46 560317 -34 560351
rect 34 560317 46 560351
rect -46 560311 46 560317
rect -46 560243 46 560249
rect -46 560209 -34 560243
rect 34 560209 46 560243
rect -46 560203 46 560209
rect -102 560159 -56 560171
rect -102 559183 -96 560159
rect -62 559183 -56 560159
rect -102 559171 -56 559183
rect 56 560159 102 560171
rect 56 559183 62 560159
rect 96 559183 102 560159
rect 56 559171 102 559183
rect -46 559133 46 559139
rect -46 559099 -34 559133
rect 34 559099 46 559133
rect -46 559093 46 559099
rect -46 559025 46 559031
rect -46 558991 -34 559025
rect 34 558991 46 559025
rect -46 558985 46 558991
rect -102 558941 -56 558953
rect -102 557965 -96 558941
rect -62 557965 -56 558941
rect -102 557953 -56 557965
rect 56 558941 102 558953
rect 56 557965 62 558941
rect 96 557965 102 558941
rect 56 557953 102 557965
rect -46 557915 46 557921
rect -46 557881 -34 557915
rect 34 557881 46 557915
rect -46 557875 46 557881
rect -46 557807 46 557813
rect -46 557773 -34 557807
rect 34 557773 46 557807
rect -46 557767 46 557773
rect -102 557723 -56 557735
rect -102 556747 -96 557723
rect -62 556747 -56 557723
rect -102 556735 -56 556747
rect 56 557723 102 557735
rect 56 556747 62 557723
rect 96 556747 102 557723
rect 56 556735 102 556747
rect -46 556697 46 556703
rect -46 556663 -34 556697
rect 34 556663 46 556697
rect -46 556657 46 556663
rect -46 556589 46 556595
rect -46 556555 -34 556589
rect 34 556555 46 556589
rect -46 556549 46 556555
rect -102 556505 -56 556517
rect -102 555529 -96 556505
rect -62 555529 -56 556505
rect -102 555517 -56 555529
rect 56 556505 102 556517
rect 56 555529 62 556505
rect 96 555529 102 556505
rect 56 555517 102 555529
rect -46 555479 46 555485
rect -46 555445 -34 555479
rect 34 555445 46 555479
rect -46 555439 46 555445
rect -46 555371 46 555377
rect -46 555337 -34 555371
rect 34 555337 46 555371
rect -46 555331 46 555337
rect -102 555287 -56 555299
rect -102 554311 -96 555287
rect -62 554311 -56 555287
rect -102 554299 -56 554311
rect 56 555287 102 555299
rect 56 554311 62 555287
rect 96 554311 102 555287
rect 56 554299 102 554311
rect -46 554261 46 554267
rect -46 554227 -34 554261
rect 34 554227 46 554261
rect -46 554221 46 554227
rect -46 554153 46 554159
rect -46 554119 -34 554153
rect 34 554119 46 554153
rect -46 554113 46 554119
rect -102 554069 -56 554081
rect -102 553093 -96 554069
rect -62 553093 -56 554069
rect -102 553081 -56 553093
rect 56 554069 102 554081
rect 56 553093 62 554069
rect 96 553093 102 554069
rect 56 553081 102 553093
rect -46 553043 46 553049
rect -46 553009 -34 553043
rect 34 553009 46 553043
rect -46 553003 46 553009
rect -46 552935 46 552941
rect -46 552901 -34 552935
rect 34 552901 46 552935
rect -46 552895 46 552901
rect -102 552851 -56 552863
rect -102 551875 -96 552851
rect -62 551875 -56 552851
rect -102 551863 -56 551875
rect 56 552851 102 552863
rect 56 551875 62 552851
rect 96 551875 102 552851
rect 56 551863 102 551875
rect -46 551825 46 551831
rect -46 551791 -34 551825
rect 34 551791 46 551825
rect -46 551785 46 551791
rect -46 551717 46 551723
rect -46 551683 -34 551717
rect 34 551683 46 551717
rect -46 551677 46 551683
rect -102 551633 -56 551645
rect -102 550657 -96 551633
rect -62 550657 -56 551633
rect -102 550645 -56 550657
rect 56 551633 102 551645
rect 56 550657 62 551633
rect 96 550657 102 551633
rect 56 550645 102 550657
rect -46 550607 46 550613
rect -46 550573 -34 550607
rect 34 550573 46 550607
rect -46 550567 46 550573
rect -46 550499 46 550505
rect -46 550465 -34 550499
rect 34 550465 46 550499
rect -46 550459 46 550465
rect -102 550415 -56 550427
rect -102 549439 -96 550415
rect -62 549439 -56 550415
rect -102 549427 -56 549439
rect 56 550415 102 550427
rect 56 549439 62 550415
rect 96 549439 102 550415
rect 56 549427 102 549439
rect -46 549389 46 549395
rect -46 549355 -34 549389
rect 34 549355 46 549389
rect -46 549349 46 549355
rect -46 549281 46 549287
rect -46 549247 -34 549281
rect 34 549247 46 549281
rect -46 549241 46 549247
rect -102 549197 -56 549209
rect -102 548221 -96 549197
rect -62 548221 -56 549197
rect -102 548209 -56 548221
rect 56 549197 102 549209
rect 56 548221 62 549197
rect 96 548221 102 549197
rect 56 548209 102 548221
rect -46 548171 46 548177
rect -46 548137 -34 548171
rect 34 548137 46 548171
rect -46 548131 46 548137
rect -46 548063 46 548069
rect -46 548029 -34 548063
rect 34 548029 46 548063
rect -46 548023 46 548029
rect -102 547979 -56 547991
rect -102 547003 -96 547979
rect -62 547003 -56 547979
rect -102 546991 -56 547003
rect 56 547979 102 547991
rect 56 547003 62 547979
rect 96 547003 102 547979
rect 56 546991 102 547003
rect -46 546953 46 546959
rect -46 546919 -34 546953
rect 34 546919 46 546953
rect -46 546913 46 546919
rect -46 546845 46 546851
rect -46 546811 -34 546845
rect 34 546811 46 546845
rect -46 546805 46 546811
rect -102 546761 -56 546773
rect -102 545785 -96 546761
rect -62 545785 -56 546761
rect -102 545773 -56 545785
rect 56 546761 102 546773
rect 56 545785 62 546761
rect 96 545785 102 546761
rect 56 545773 102 545785
rect -46 545735 46 545741
rect -46 545701 -34 545735
rect 34 545701 46 545735
rect -46 545695 46 545701
rect -46 545627 46 545633
rect -46 545593 -34 545627
rect 34 545593 46 545627
rect -46 545587 46 545593
rect -102 545543 -56 545555
rect -102 544567 -96 545543
rect -62 544567 -56 545543
rect -102 544555 -56 544567
rect 56 545543 102 545555
rect 56 544567 62 545543
rect 96 544567 102 545543
rect 56 544555 102 544567
rect -46 544517 46 544523
rect -46 544483 -34 544517
rect 34 544483 46 544517
rect -46 544477 46 544483
rect -46 544409 46 544415
rect -46 544375 -34 544409
rect 34 544375 46 544409
rect -46 544369 46 544375
rect -102 544325 -56 544337
rect -102 543349 -96 544325
rect -62 543349 -56 544325
rect -102 543337 -56 543349
rect 56 544325 102 544337
rect 56 543349 62 544325
rect 96 543349 102 544325
rect 56 543337 102 543349
rect -46 543299 46 543305
rect -46 543265 -34 543299
rect 34 543265 46 543299
rect -46 543259 46 543265
rect -46 543191 46 543197
rect -46 543157 -34 543191
rect 34 543157 46 543191
rect -46 543151 46 543157
rect -102 543107 -56 543119
rect -102 542131 -96 543107
rect -62 542131 -56 543107
rect -102 542119 -56 542131
rect 56 543107 102 543119
rect 56 542131 62 543107
rect 96 542131 102 543107
rect 56 542119 102 542131
rect -46 542081 46 542087
rect -46 542047 -34 542081
rect 34 542047 46 542081
rect -46 542041 46 542047
rect -46 541973 46 541979
rect -46 541939 -34 541973
rect 34 541939 46 541973
rect -46 541933 46 541939
rect -102 541889 -56 541901
rect -102 540913 -96 541889
rect -62 540913 -56 541889
rect -102 540901 -56 540913
rect 56 541889 102 541901
rect 56 540913 62 541889
rect 96 540913 102 541889
rect 56 540901 102 540913
rect -46 540863 46 540869
rect -46 540829 -34 540863
rect 34 540829 46 540863
rect -46 540823 46 540829
rect -46 540755 46 540761
rect -46 540721 -34 540755
rect 34 540721 46 540755
rect -46 540715 46 540721
rect -102 540671 -56 540683
rect -102 539695 -96 540671
rect -62 539695 -56 540671
rect -102 539683 -56 539695
rect 56 540671 102 540683
rect 56 539695 62 540671
rect 96 539695 102 540671
rect 56 539683 102 539695
rect -46 539645 46 539651
rect -46 539611 -34 539645
rect 34 539611 46 539645
rect -46 539605 46 539611
rect -46 539537 46 539543
rect -46 539503 -34 539537
rect 34 539503 46 539537
rect -46 539497 46 539503
rect -102 539453 -56 539465
rect -102 538477 -96 539453
rect -62 538477 -56 539453
rect -102 538465 -56 538477
rect 56 539453 102 539465
rect 56 538477 62 539453
rect 96 538477 102 539453
rect 56 538465 102 538477
rect -46 538427 46 538433
rect -46 538393 -34 538427
rect 34 538393 46 538427
rect -46 538387 46 538393
rect -46 538319 46 538325
rect -46 538285 -34 538319
rect 34 538285 46 538319
rect -46 538279 46 538285
rect -102 538235 -56 538247
rect -102 537259 -96 538235
rect -62 537259 -56 538235
rect -102 537247 -56 537259
rect 56 538235 102 538247
rect 56 537259 62 538235
rect 96 537259 102 538235
rect 56 537247 102 537259
rect -46 537209 46 537215
rect -46 537175 -34 537209
rect 34 537175 46 537209
rect -46 537169 46 537175
rect -46 537101 46 537107
rect -46 537067 -34 537101
rect 34 537067 46 537101
rect -46 537061 46 537067
rect -102 537017 -56 537029
rect -102 536041 -96 537017
rect -62 536041 -56 537017
rect -102 536029 -56 536041
rect 56 537017 102 537029
rect 56 536041 62 537017
rect 96 536041 102 537017
rect 56 536029 102 536041
rect -46 535991 46 535997
rect -46 535957 -34 535991
rect 34 535957 46 535991
rect -46 535951 46 535957
rect -46 535883 46 535889
rect -46 535849 -34 535883
rect 34 535849 46 535883
rect -46 535843 46 535849
rect -102 535799 -56 535811
rect -102 534823 -96 535799
rect -62 534823 -56 535799
rect -102 534811 -56 534823
rect 56 535799 102 535811
rect 56 534823 62 535799
rect 96 534823 102 535799
rect 56 534811 102 534823
rect -46 534773 46 534779
rect -46 534739 -34 534773
rect 34 534739 46 534773
rect -46 534733 46 534739
rect -46 534665 46 534671
rect -46 534631 -34 534665
rect 34 534631 46 534665
rect -46 534625 46 534631
rect -102 534581 -56 534593
rect -102 533605 -96 534581
rect -62 533605 -56 534581
rect -102 533593 -56 533605
rect 56 534581 102 534593
rect 56 533605 62 534581
rect 96 533605 102 534581
rect 56 533593 102 533605
rect -46 533555 46 533561
rect -46 533521 -34 533555
rect 34 533521 46 533555
rect -46 533515 46 533521
rect -46 533447 46 533453
rect -46 533413 -34 533447
rect 34 533413 46 533447
rect -46 533407 46 533413
rect -102 533363 -56 533375
rect -102 532387 -96 533363
rect -62 532387 -56 533363
rect -102 532375 -56 532387
rect 56 533363 102 533375
rect 56 532387 62 533363
rect 96 532387 102 533363
rect 56 532375 102 532387
rect -46 532337 46 532343
rect -46 532303 -34 532337
rect 34 532303 46 532337
rect -46 532297 46 532303
rect -46 532229 46 532235
rect -46 532195 -34 532229
rect 34 532195 46 532229
rect -46 532189 46 532195
rect -102 532145 -56 532157
rect -102 531169 -96 532145
rect -62 531169 -56 532145
rect -102 531157 -56 531169
rect 56 532145 102 532157
rect 56 531169 62 532145
rect 96 531169 102 532145
rect 56 531157 102 531169
rect -46 531119 46 531125
rect -46 531085 -34 531119
rect 34 531085 46 531119
rect -46 531079 46 531085
rect -46 531011 46 531017
rect -46 530977 -34 531011
rect 34 530977 46 531011
rect -46 530971 46 530977
rect -102 530927 -56 530939
rect -102 529951 -96 530927
rect -62 529951 -56 530927
rect -102 529939 -56 529951
rect 56 530927 102 530939
rect 56 529951 62 530927
rect 96 529951 102 530927
rect 56 529939 102 529951
rect -46 529901 46 529907
rect -46 529867 -34 529901
rect 34 529867 46 529901
rect -46 529861 46 529867
rect -46 529793 46 529799
rect -46 529759 -34 529793
rect 34 529759 46 529793
rect -46 529753 46 529759
rect -102 529709 -56 529721
rect -102 528733 -96 529709
rect -62 528733 -56 529709
rect -102 528721 -56 528733
rect 56 529709 102 529721
rect 56 528733 62 529709
rect 96 528733 102 529709
rect 56 528721 102 528733
rect -46 528683 46 528689
rect -46 528649 -34 528683
rect 34 528649 46 528683
rect -46 528643 46 528649
rect -46 528575 46 528581
rect -46 528541 -34 528575
rect 34 528541 46 528575
rect -46 528535 46 528541
rect -102 528491 -56 528503
rect -102 527515 -96 528491
rect -62 527515 -56 528491
rect -102 527503 -56 527515
rect 56 528491 102 528503
rect 56 527515 62 528491
rect 96 527515 102 528491
rect 56 527503 102 527515
rect -46 527465 46 527471
rect -46 527431 -34 527465
rect 34 527431 46 527465
rect -46 527425 46 527431
rect -46 527357 46 527363
rect -46 527323 -34 527357
rect 34 527323 46 527357
rect -46 527317 46 527323
rect -102 527273 -56 527285
rect -102 526297 -96 527273
rect -62 526297 -56 527273
rect -102 526285 -56 526297
rect 56 527273 102 527285
rect 56 526297 62 527273
rect 96 526297 102 527273
rect 56 526285 102 526297
rect -46 526247 46 526253
rect -46 526213 -34 526247
rect 34 526213 46 526247
rect -46 526207 46 526213
rect -46 526139 46 526145
rect -46 526105 -34 526139
rect 34 526105 46 526139
rect -46 526099 46 526105
rect -102 526055 -56 526067
rect -102 525079 -96 526055
rect -62 525079 -56 526055
rect -102 525067 -56 525079
rect 56 526055 102 526067
rect 56 525079 62 526055
rect 96 525079 102 526055
rect 56 525067 102 525079
rect -46 525029 46 525035
rect -46 524995 -34 525029
rect 34 524995 46 525029
rect -46 524989 46 524995
rect -46 524921 46 524927
rect -46 524887 -34 524921
rect 34 524887 46 524921
rect -46 524881 46 524887
rect -102 524837 -56 524849
rect -102 523861 -96 524837
rect -62 523861 -56 524837
rect -102 523849 -56 523861
rect 56 524837 102 524849
rect 56 523861 62 524837
rect 96 523861 102 524837
rect 56 523849 102 523861
rect -46 523811 46 523817
rect -46 523777 -34 523811
rect 34 523777 46 523811
rect -46 523771 46 523777
rect -46 523703 46 523709
rect -46 523669 -34 523703
rect 34 523669 46 523703
rect -46 523663 46 523669
rect -102 523619 -56 523631
rect -102 522643 -96 523619
rect -62 522643 -56 523619
rect -102 522631 -56 522643
rect 56 523619 102 523631
rect 56 522643 62 523619
rect 96 522643 102 523619
rect 56 522631 102 522643
rect -46 522593 46 522599
rect -46 522559 -34 522593
rect 34 522559 46 522593
rect -46 522553 46 522559
rect -46 522485 46 522491
rect -46 522451 -34 522485
rect 34 522451 46 522485
rect -46 522445 46 522451
rect -102 522401 -56 522413
rect -102 521425 -96 522401
rect -62 521425 -56 522401
rect -102 521413 -56 521425
rect 56 522401 102 522413
rect 56 521425 62 522401
rect 96 521425 102 522401
rect 56 521413 102 521425
rect -46 521375 46 521381
rect -46 521341 -34 521375
rect 34 521341 46 521375
rect -46 521335 46 521341
rect -46 521267 46 521273
rect -46 521233 -34 521267
rect 34 521233 46 521267
rect -46 521227 46 521233
rect -102 521183 -56 521195
rect -102 520207 -96 521183
rect -62 520207 -56 521183
rect -102 520195 -56 520207
rect 56 521183 102 521195
rect 56 520207 62 521183
rect 96 520207 102 521183
rect 56 520195 102 520207
rect -46 520157 46 520163
rect -46 520123 -34 520157
rect 34 520123 46 520157
rect -46 520117 46 520123
rect -46 520049 46 520055
rect -46 520015 -34 520049
rect 34 520015 46 520049
rect -46 520009 46 520015
rect -102 519965 -56 519977
rect -102 518989 -96 519965
rect -62 518989 -56 519965
rect -102 518977 -56 518989
rect 56 519965 102 519977
rect 56 518989 62 519965
rect 96 518989 102 519965
rect 56 518977 102 518989
rect -46 518939 46 518945
rect -46 518905 -34 518939
rect 34 518905 46 518939
rect -46 518899 46 518905
rect -46 518831 46 518837
rect -46 518797 -34 518831
rect 34 518797 46 518831
rect -46 518791 46 518797
rect -102 518747 -56 518759
rect -102 517771 -96 518747
rect -62 517771 -56 518747
rect -102 517759 -56 517771
rect 56 518747 102 518759
rect 56 517771 62 518747
rect 96 517771 102 518747
rect 56 517759 102 517771
rect -46 517721 46 517727
rect -46 517687 -34 517721
rect 34 517687 46 517721
rect -46 517681 46 517687
rect -46 517613 46 517619
rect -46 517579 -34 517613
rect 34 517579 46 517613
rect -46 517573 46 517579
rect -102 517529 -56 517541
rect -102 516553 -96 517529
rect -62 516553 -56 517529
rect -102 516541 -56 516553
rect 56 517529 102 517541
rect 56 516553 62 517529
rect 96 516553 102 517529
rect 56 516541 102 516553
rect -46 516503 46 516509
rect -46 516469 -34 516503
rect 34 516469 46 516503
rect -46 516463 46 516469
rect -46 516395 46 516401
rect -46 516361 -34 516395
rect 34 516361 46 516395
rect -46 516355 46 516361
rect -102 516311 -56 516323
rect -102 515335 -96 516311
rect -62 515335 -56 516311
rect -102 515323 -56 515335
rect 56 516311 102 516323
rect 56 515335 62 516311
rect 96 515335 102 516311
rect 56 515323 102 515335
rect -46 515285 46 515291
rect -46 515251 -34 515285
rect 34 515251 46 515285
rect -46 515245 46 515251
rect -46 515177 46 515183
rect -46 515143 -34 515177
rect 34 515143 46 515177
rect -46 515137 46 515143
rect -102 515093 -56 515105
rect -102 514117 -96 515093
rect -62 514117 -56 515093
rect -102 514105 -56 514117
rect 56 515093 102 515105
rect 56 514117 62 515093
rect 96 514117 102 515093
rect 56 514105 102 514117
rect -46 514067 46 514073
rect -46 514033 -34 514067
rect 34 514033 46 514067
rect -46 514027 46 514033
rect -46 513959 46 513965
rect -46 513925 -34 513959
rect 34 513925 46 513959
rect -46 513919 46 513925
rect -102 513875 -56 513887
rect -102 512899 -96 513875
rect -62 512899 -56 513875
rect -102 512887 -56 512899
rect 56 513875 102 513887
rect 56 512899 62 513875
rect 96 512899 102 513875
rect 56 512887 102 512899
rect -46 512849 46 512855
rect -46 512815 -34 512849
rect 34 512815 46 512849
rect -46 512809 46 512815
rect -46 512741 46 512747
rect -46 512707 -34 512741
rect 34 512707 46 512741
rect -46 512701 46 512707
rect -102 512657 -56 512669
rect -102 511681 -96 512657
rect -62 511681 -56 512657
rect -102 511669 -56 511681
rect 56 512657 102 512669
rect 56 511681 62 512657
rect 96 511681 102 512657
rect 56 511669 102 511681
rect -46 511631 46 511637
rect -46 511597 -34 511631
rect 34 511597 46 511631
rect -46 511591 46 511597
rect -46 511523 46 511529
rect -46 511489 -34 511523
rect 34 511489 46 511523
rect -46 511483 46 511489
rect -102 511439 -56 511451
rect -102 510463 -96 511439
rect -62 510463 -56 511439
rect -102 510451 -56 510463
rect 56 511439 102 511451
rect 56 510463 62 511439
rect 96 510463 102 511439
rect 56 510451 102 510463
rect -46 510413 46 510419
rect -46 510379 -34 510413
rect 34 510379 46 510413
rect -46 510373 46 510379
rect -46 510305 46 510311
rect -46 510271 -34 510305
rect 34 510271 46 510305
rect -46 510265 46 510271
rect -102 510221 -56 510233
rect -102 509245 -96 510221
rect -62 509245 -56 510221
rect -102 509233 -56 509245
rect 56 510221 102 510233
rect 56 509245 62 510221
rect 96 509245 102 510221
rect 56 509233 102 509245
rect -46 509195 46 509201
rect -46 509161 -34 509195
rect 34 509161 46 509195
rect -46 509155 46 509161
rect -46 509087 46 509093
rect -46 509053 -34 509087
rect 34 509053 46 509087
rect -46 509047 46 509053
rect -102 509003 -56 509015
rect -102 508027 -96 509003
rect -62 508027 -56 509003
rect -102 508015 -56 508027
rect 56 509003 102 509015
rect 56 508027 62 509003
rect 96 508027 102 509003
rect 56 508015 102 508027
rect -46 507977 46 507983
rect -46 507943 -34 507977
rect 34 507943 46 507977
rect -46 507937 46 507943
rect -46 507869 46 507875
rect -46 507835 -34 507869
rect 34 507835 46 507869
rect -46 507829 46 507835
rect -102 507785 -56 507797
rect -102 506809 -96 507785
rect -62 506809 -56 507785
rect -102 506797 -56 506809
rect 56 507785 102 507797
rect 56 506809 62 507785
rect 96 506809 102 507785
rect 56 506797 102 506809
rect -46 506759 46 506765
rect -46 506725 -34 506759
rect 34 506725 46 506759
rect -46 506719 46 506725
rect -46 506651 46 506657
rect -46 506617 -34 506651
rect 34 506617 46 506651
rect -46 506611 46 506617
rect -102 506567 -56 506579
rect -102 505591 -96 506567
rect -62 505591 -56 506567
rect -102 505579 -56 505591
rect 56 506567 102 506579
rect 56 505591 62 506567
rect 96 505591 102 506567
rect 56 505579 102 505591
rect -46 505541 46 505547
rect -46 505507 -34 505541
rect 34 505507 46 505541
rect -46 505501 46 505507
rect -46 505433 46 505439
rect -46 505399 -34 505433
rect 34 505399 46 505433
rect -46 505393 46 505399
rect -102 505349 -56 505361
rect -102 504373 -96 505349
rect -62 504373 -56 505349
rect -102 504361 -56 504373
rect 56 505349 102 505361
rect 56 504373 62 505349
rect 96 504373 102 505349
rect 56 504361 102 504373
rect -46 504323 46 504329
rect -46 504289 -34 504323
rect 34 504289 46 504323
rect -46 504283 46 504289
rect -46 504215 46 504221
rect -46 504181 -34 504215
rect 34 504181 46 504215
rect -46 504175 46 504181
rect -102 504131 -56 504143
rect -102 503155 -96 504131
rect -62 503155 -56 504131
rect -102 503143 -56 503155
rect 56 504131 102 504143
rect 56 503155 62 504131
rect 96 503155 102 504131
rect 56 503143 102 503155
rect -46 503105 46 503111
rect -46 503071 -34 503105
rect 34 503071 46 503105
rect -46 503065 46 503071
rect -46 502997 46 503003
rect -46 502963 -34 502997
rect 34 502963 46 502997
rect -46 502957 46 502963
rect -102 502913 -56 502925
rect -102 501937 -96 502913
rect -62 501937 -56 502913
rect -102 501925 -56 501937
rect 56 502913 102 502925
rect 56 501937 62 502913
rect 96 501937 102 502913
rect 56 501925 102 501937
rect -46 501887 46 501893
rect -46 501853 -34 501887
rect 34 501853 46 501887
rect -46 501847 46 501853
rect -46 501779 46 501785
rect -46 501745 -34 501779
rect 34 501745 46 501779
rect -46 501739 46 501745
rect -102 501695 -56 501707
rect -102 500719 -96 501695
rect -62 500719 -56 501695
rect -102 500707 -56 500719
rect 56 501695 102 501707
rect 56 500719 62 501695
rect 96 500719 102 501695
rect 56 500707 102 500719
rect -46 500669 46 500675
rect -46 500635 -34 500669
rect 34 500635 46 500669
rect -46 500629 46 500635
rect -46 500561 46 500567
rect -46 500527 -34 500561
rect 34 500527 46 500561
rect -46 500521 46 500527
rect -102 500477 -56 500489
rect -102 499501 -96 500477
rect -62 499501 -56 500477
rect -102 499489 -56 499501
rect 56 500477 102 500489
rect 56 499501 62 500477
rect 96 499501 102 500477
rect 56 499489 102 499501
rect -46 499451 46 499457
rect -46 499417 -34 499451
rect 34 499417 46 499451
rect -46 499411 46 499417
rect -46 499343 46 499349
rect -46 499309 -34 499343
rect 34 499309 46 499343
rect -46 499303 46 499309
rect -102 499259 -56 499271
rect -102 498283 -96 499259
rect -62 498283 -56 499259
rect -102 498271 -56 498283
rect 56 499259 102 499271
rect 56 498283 62 499259
rect 96 498283 102 499259
rect 56 498271 102 498283
rect -46 498233 46 498239
rect -46 498199 -34 498233
rect 34 498199 46 498233
rect -46 498193 46 498199
rect -46 498125 46 498131
rect -46 498091 -34 498125
rect 34 498091 46 498125
rect -46 498085 46 498091
rect -102 498041 -56 498053
rect -102 497065 -96 498041
rect -62 497065 -56 498041
rect -102 497053 -56 497065
rect 56 498041 102 498053
rect 56 497065 62 498041
rect 96 497065 102 498041
rect 56 497053 102 497065
rect -46 497015 46 497021
rect -46 496981 -34 497015
rect 34 496981 46 497015
rect -46 496975 46 496981
rect -46 496907 46 496913
rect -46 496873 -34 496907
rect 34 496873 46 496907
rect -46 496867 46 496873
rect -102 496823 -56 496835
rect -102 495847 -96 496823
rect -62 495847 -56 496823
rect -102 495835 -56 495847
rect 56 496823 102 496835
rect 56 495847 62 496823
rect 96 495847 102 496823
rect 56 495835 102 495847
rect -46 495797 46 495803
rect -46 495763 -34 495797
rect 34 495763 46 495797
rect -46 495757 46 495763
rect -46 495689 46 495695
rect -46 495655 -34 495689
rect 34 495655 46 495689
rect -46 495649 46 495655
rect -102 495605 -56 495617
rect -102 494629 -96 495605
rect -62 494629 -56 495605
rect -102 494617 -56 494629
rect 56 495605 102 495617
rect 56 494629 62 495605
rect 96 494629 102 495605
rect 56 494617 102 494629
rect -46 494579 46 494585
rect -46 494545 -34 494579
rect 34 494545 46 494579
rect -46 494539 46 494545
rect -46 494471 46 494477
rect -46 494437 -34 494471
rect 34 494437 46 494471
rect -46 494431 46 494437
rect -102 494387 -56 494399
rect -102 493411 -96 494387
rect -62 493411 -56 494387
rect -102 493399 -56 493411
rect 56 494387 102 494399
rect 56 493411 62 494387
rect 96 493411 102 494387
rect 56 493399 102 493411
rect -46 493361 46 493367
rect -46 493327 -34 493361
rect 34 493327 46 493361
rect -46 493321 46 493327
rect -46 493253 46 493259
rect -46 493219 -34 493253
rect 34 493219 46 493253
rect -46 493213 46 493219
rect -102 493169 -56 493181
rect -102 492193 -96 493169
rect -62 492193 -56 493169
rect -102 492181 -56 492193
rect 56 493169 102 493181
rect 56 492193 62 493169
rect 96 492193 102 493169
rect 56 492181 102 492193
rect -46 492143 46 492149
rect -46 492109 -34 492143
rect 34 492109 46 492143
rect -46 492103 46 492109
rect -46 492035 46 492041
rect -46 492001 -34 492035
rect 34 492001 46 492035
rect -46 491995 46 492001
rect -102 491951 -56 491963
rect -102 490975 -96 491951
rect -62 490975 -56 491951
rect -102 490963 -56 490975
rect 56 491951 102 491963
rect 56 490975 62 491951
rect 96 490975 102 491951
rect 56 490963 102 490975
rect -46 490925 46 490931
rect -46 490891 -34 490925
rect 34 490891 46 490925
rect -46 490885 46 490891
rect -46 490817 46 490823
rect -46 490783 -34 490817
rect 34 490783 46 490817
rect -46 490777 46 490783
rect -102 490733 -56 490745
rect -102 489757 -96 490733
rect -62 489757 -56 490733
rect -102 489745 -56 489757
rect 56 490733 102 490745
rect 56 489757 62 490733
rect 96 489757 102 490733
rect 56 489745 102 489757
rect -46 489707 46 489713
rect -46 489673 -34 489707
rect 34 489673 46 489707
rect -46 489667 46 489673
rect -46 489599 46 489605
rect -46 489565 -34 489599
rect 34 489565 46 489599
rect -46 489559 46 489565
rect -102 489515 -56 489527
rect -102 488539 -96 489515
rect -62 488539 -56 489515
rect -102 488527 -56 488539
rect 56 489515 102 489527
rect 56 488539 62 489515
rect 96 488539 102 489515
rect 56 488527 102 488539
rect -46 488489 46 488495
rect -46 488455 -34 488489
rect 34 488455 46 488489
rect -46 488449 46 488455
rect -46 488381 46 488387
rect -46 488347 -34 488381
rect 34 488347 46 488381
rect -46 488341 46 488347
rect -102 488297 -56 488309
rect -102 487321 -96 488297
rect -62 487321 -56 488297
rect -102 487309 -56 487321
rect 56 488297 102 488309
rect 56 487321 62 488297
rect 96 487321 102 488297
rect 56 487309 102 487321
rect -46 487271 46 487277
rect -46 487237 -34 487271
rect 34 487237 46 487271
rect -46 487231 46 487237
rect -46 487163 46 487169
rect -46 487129 -34 487163
rect 34 487129 46 487163
rect -46 487123 46 487129
rect -102 487079 -56 487091
rect -102 486103 -96 487079
rect -62 486103 -56 487079
rect -102 486091 -56 486103
rect 56 487079 102 487091
rect 56 486103 62 487079
rect 96 486103 102 487079
rect 56 486091 102 486103
rect -46 486053 46 486059
rect -46 486019 -34 486053
rect 34 486019 46 486053
rect -46 486013 46 486019
rect -46 485945 46 485951
rect -46 485911 -34 485945
rect 34 485911 46 485945
rect -46 485905 46 485911
rect -102 485861 -56 485873
rect -102 484885 -96 485861
rect -62 484885 -56 485861
rect -102 484873 -56 484885
rect 56 485861 102 485873
rect 56 484885 62 485861
rect 96 484885 102 485861
rect 56 484873 102 484885
rect -46 484835 46 484841
rect -46 484801 -34 484835
rect 34 484801 46 484835
rect -46 484795 46 484801
rect -46 484727 46 484733
rect -46 484693 -34 484727
rect 34 484693 46 484727
rect -46 484687 46 484693
rect -102 484643 -56 484655
rect -102 483667 -96 484643
rect -62 483667 -56 484643
rect -102 483655 -56 483667
rect 56 484643 102 484655
rect 56 483667 62 484643
rect 96 483667 102 484643
rect 56 483655 102 483667
rect -46 483617 46 483623
rect -46 483583 -34 483617
rect 34 483583 46 483617
rect -46 483577 46 483583
rect -46 483509 46 483515
rect -46 483475 -34 483509
rect 34 483475 46 483509
rect -46 483469 46 483475
rect -102 483425 -56 483437
rect -102 482449 -96 483425
rect -62 482449 -56 483425
rect -102 482437 -56 482449
rect 56 483425 102 483437
rect 56 482449 62 483425
rect 96 482449 102 483425
rect 56 482437 102 482449
rect -46 482399 46 482405
rect -46 482365 -34 482399
rect 34 482365 46 482399
rect -46 482359 46 482365
rect -46 482291 46 482297
rect -46 482257 -34 482291
rect 34 482257 46 482291
rect -46 482251 46 482257
rect -102 482207 -56 482219
rect -102 481231 -96 482207
rect -62 481231 -56 482207
rect -102 481219 -56 481231
rect 56 482207 102 482219
rect 56 481231 62 482207
rect 96 481231 102 482207
rect 56 481219 102 481231
rect -46 481181 46 481187
rect -46 481147 -34 481181
rect 34 481147 46 481181
rect -46 481141 46 481147
rect -46 481073 46 481079
rect -46 481039 -34 481073
rect 34 481039 46 481073
rect -46 481033 46 481039
rect -102 480989 -56 481001
rect -102 480013 -96 480989
rect -62 480013 -56 480989
rect -102 480001 -56 480013
rect 56 480989 102 481001
rect 56 480013 62 480989
rect 96 480013 102 480989
rect 56 480001 102 480013
rect -46 479963 46 479969
rect -46 479929 -34 479963
rect 34 479929 46 479963
rect -46 479923 46 479929
rect -46 479855 46 479861
rect -46 479821 -34 479855
rect 34 479821 46 479855
rect -46 479815 46 479821
rect -102 479771 -56 479783
rect -102 478795 -96 479771
rect -62 478795 -56 479771
rect -102 478783 -56 478795
rect 56 479771 102 479783
rect 56 478795 62 479771
rect 96 478795 102 479771
rect 56 478783 102 478795
rect -46 478745 46 478751
rect -46 478711 -34 478745
rect 34 478711 46 478745
rect -46 478705 46 478711
rect -46 478637 46 478643
rect -46 478603 -34 478637
rect 34 478603 46 478637
rect -46 478597 46 478603
rect -102 478553 -56 478565
rect -102 477577 -96 478553
rect -62 477577 -56 478553
rect -102 477565 -56 477577
rect 56 478553 102 478565
rect 56 477577 62 478553
rect 96 477577 102 478553
rect 56 477565 102 477577
rect -46 477527 46 477533
rect -46 477493 -34 477527
rect 34 477493 46 477527
rect -46 477487 46 477493
rect -46 477419 46 477425
rect -46 477385 -34 477419
rect 34 477385 46 477419
rect -46 477379 46 477385
rect -102 477335 -56 477347
rect -102 476359 -96 477335
rect -62 476359 -56 477335
rect -102 476347 -56 476359
rect 56 477335 102 477347
rect 56 476359 62 477335
rect 96 476359 102 477335
rect 56 476347 102 476359
rect -46 476309 46 476315
rect -46 476275 -34 476309
rect 34 476275 46 476309
rect -46 476269 46 476275
rect -46 476201 46 476207
rect -46 476167 -34 476201
rect 34 476167 46 476201
rect -46 476161 46 476167
rect -102 476117 -56 476129
rect -102 475141 -96 476117
rect -62 475141 -56 476117
rect -102 475129 -56 475141
rect 56 476117 102 476129
rect 56 475141 62 476117
rect 96 475141 102 476117
rect 56 475129 102 475141
rect -46 475091 46 475097
rect -46 475057 -34 475091
rect 34 475057 46 475091
rect -46 475051 46 475057
rect -46 474983 46 474989
rect -46 474949 -34 474983
rect 34 474949 46 474983
rect -46 474943 46 474949
rect -102 474899 -56 474911
rect -102 473923 -96 474899
rect -62 473923 -56 474899
rect -102 473911 -56 473923
rect 56 474899 102 474911
rect 56 473923 62 474899
rect 96 473923 102 474899
rect 56 473911 102 473923
rect -46 473873 46 473879
rect -46 473839 -34 473873
rect 34 473839 46 473873
rect -46 473833 46 473839
rect -46 473765 46 473771
rect -46 473731 -34 473765
rect 34 473731 46 473765
rect -46 473725 46 473731
rect -102 473681 -56 473693
rect -102 472705 -96 473681
rect -62 472705 -56 473681
rect -102 472693 -56 472705
rect 56 473681 102 473693
rect 56 472705 62 473681
rect 96 472705 102 473681
rect 56 472693 102 472705
rect -46 472655 46 472661
rect -46 472621 -34 472655
rect 34 472621 46 472655
rect -46 472615 46 472621
rect -46 472547 46 472553
rect -46 472513 -34 472547
rect 34 472513 46 472547
rect -46 472507 46 472513
rect -102 472463 -56 472475
rect -102 471487 -96 472463
rect -62 471487 -56 472463
rect -102 471475 -56 471487
rect 56 472463 102 472475
rect 56 471487 62 472463
rect 96 471487 102 472463
rect 56 471475 102 471487
rect -46 471437 46 471443
rect -46 471403 -34 471437
rect 34 471403 46 471437
rect -46 471397 46 471403
rect -46 471329 46 471335
rect -46 471295 -34 471329
rect 34 471295 46 471329
rect -46 471289 46 471295
rect -102 471245 -56 471257
rect -102 470269 -96 471245
rect -62 470269 -56 471245
rect -102 470257 -56 470269
rect 56 471245 102 471257
rect 56 470269 62 471245
rect 96 470269 102 471245
rect 56 470257 102 470269
rect -46 470219 46 470225
rect -46 470185 -34 470219
rect 34 470185 46 470219
rect -46 470179 46 470185
rect -46 470111 46 470117
rect -46 470077 -34 470111
rect 34 470077 46 470111
rect -46 470071 46 470077
rect -102 470027 -56 470039
rect -102 469051 -96 470027
rect -62 469051 -56 470027
rect -102 469039 -56 469051
rect 56 470027 102 470039
rect 56 469051 62 470027
rect 96 469051 102 470027
rect 56 469039 102 469051
rect -46 469001 46 469007
rect -46 468967 -34 469001
rect 34 468967 46 469001
rect -46 468961 46 468967
rect -46 468893 46 468899
rect -46 468859 -34 468893
rect 34 468859 46 468893
rect -46 468853 46 468859
rect -102 468809 -56 468821
rect -102 467833 -96 468809
rect -62 467833 -56 468809
rect -102 467821 -56 467833
rect 56 468809 102 468821
rect 56 467833 62 468809
rect 96 467833 102 468809
rect 56 467821 102 467833
rect -46 467783 46 467789
rect -46 467749 -34 467783
rect 34 467749 46 467783
rect -46 467743 46 467749
rect -46 467675 46 467681
rect -46 467641 -34 467675
rect 34 467641 46 467675
rect -46 467635 46 467641
rect -102 467591 -56 467603
rect -102 466615 -96 467591
rect -62 466615 -56 467591
rect -102 466603 -56 466615
rect 56 467591 102 467603
rect 56 466615 62 467591
rect 96 466615 102 467591
rect 56 466603 102 466615
rect -46 466565 46 466571
rect -46 466531 -34 466565
rect 34 466531 46 466565
rect -46 466525 46 466531
rect -46 466457 46 466463
rect -46 466423 -34 466457
rect 34 466423 46 466457
rect -46 466417 46 466423
rect -102 466373 -56 466385
rect -102 465397 -96 466373
rect -62 465397 -56 466373
rect -102 465385 -56 465397
rect 56 466373 102 466385
rect 56 465397 62 466373
rect 96 465397 102 466373
rect 56 465385 102 465397
rect -46 465347 46 465353
rect -46 465313 -34 465347
rect 34 465313 46 465347
rect -46 465307 46 465313
rect -46 465239 46 465245
rect -46 465205 -34 465239
rect 34 465205 46 465239
rect -46 465199 46 465205
rect -102 465155 -56 465167
rect -102 464179 -96 465155
rect -62 464179 -56 465155
rect -102 464167 -56 464179
rect 56 465155 102 465167
rect 56 464179 62 465155
rect 96 464179 102 465155
rect 56 464167 102 464179
rect -46 464129 46 464135
rect -46 464095 -34 464129
rect 34 464095 46 464129
rect -46 464089 46 464095
rect -46 464021 46 464027
rect -46 463987 -34 464021
rect 34 463987 46 464021
rect -46 463981 46 463987
rect -102 463937 -56 463949
rect -102 462961 -96 463937
rect -62 462961 -56 463937
rect -102 462949 -56 462961
rect 56 463937 102 463949
rect 56 462961 62 463937
rect 96 462961 102 463937
rect 56 462949 102 462961
rect -46 462911 46 462917
rect -46 462877 -34 462911
rect 34 462877 46 462911
rect -46 462871 46 462877
rect -46 462803 46 462809
rect -46 462769 -34 462803
rect 34 462769 46 462803
rect -46 462763 46 462769
rect -102 462719 -56 462731
rect -102 461743 -96 462719
rect -62 461743 -56 462719
rect -102 461731 -56 461743
rect 56 462719 102 462731
rect 56 461743 62 462719
rect 96 461743 102 462719
rect 56 461731 102 461743
rect -46 461693 46 461699
rect -46 461659 -34 461693
rect 34 461659 46 461693
rect -46 461653 46 461659
rect -46 461585 46 461591
rect -46 461551 -34 461585
rect 34 461551 46 461585
rect -46 461545 46 461551
rect -102 461501 -56 461513
rect -102 460525 -96 461501
rect -62 460525 -56 461501
rect -102 460513 -56 460525
rect 56 461501 102 461513
rect 56 460525 62 461501
rect 96 460525 102 461501
rect 56 460513 102 460525
rect -46 460475 46 460481
rect -46 460441 -34 460475
rect 34 460441 46 460475
rect -46 460435 46 460441
rect -46 460367 46 460373
rect -46 460333 -34 460367
rect 34 460333 46 460367
rect -46 460327 46 460333
rect -102 460283 -56 460295
rect -102 459307 -96 460283
rect -62 459307 -56 460283
rect -102 459295 -56 459307
rect 56 460283 102 460295
rect 56 459307 62 460283
rect 96 459307 102 460283
rect 56 459295 102 459307
rect -46 459257 46 459263
rect -46 459223 -34 459257
rect 34 459223 46 459257
rect -46 459217 46 459223
rect -46 459149 46 459155
rect -46 459115 -34 459149
rect 34 459115 46 459149
rect -46 459109 46 459115
rect -102 459065 -56 459077
rect -102 458089 -96 459065
rect -62 458089 -56 459065
rect -102 458077 -56 458089
rect 56 459065 102 459077
rect 56 458089 62 459065
rect 96 458089 102 459065
rect 56 458077 102 458089
rect -46 458039 46 458045
rect -46 458005 -34 458039
rect 34 458005 46 458039
rect -46 457999 46 458005
rect -46 457931 46 457937
rect -46 457897 -34 457931
rect 34 457897 46 457931
rect -46 457891 46 457897
rect -102 457847 -56 457859
rect -102 456871 -96 457847
rect -62 456871 -56 457847
rect -102 456859 -56 456871
rect 56 457847 102 457859
rect 56 456871 62 457847
rect 96 456871 102 457847
rect 56 456859 102 456871
rect -46 456821 46 456827
rect -46 456787 -34 456821
rect 34 456787 46 456821
rect -46 456781 46 456787
rect -46 456713 46 456719
rect -46 456679 -34 456713
rect 34 456679 46 456713
rect -46 456673 46 456679
rect -102 456629 -56 456641
rect -102 455653 -96 456629
rect -62 455653 -56 456629
rect -102 455641 -56 455653
rect 56 456629 102 456641
rect 56 455653 62 456629
rect 96 455653 102 456629
rect 56 455641 102 455653
rect -46 455603 46 455609
rect -46 455569 -34 455603
rect 34 455569 46 455603
rect -46 455563 46 455569
rect -46 455495 46 455501
rect -46 455461 -34 455495
rect 34 455461 46 455495
rect -46 455455 46 455461
rect -102 455411 -56 455423
rect -102 454435 -96 455411
rect -62 454435 -56 455411
rect -102 454423 -56 454435
rect 56 455411 102 455423
rect 56 454435 62 455411
rect 96 454435 102 455411
rect 56 454423 102 454435
rect -46 454385 46 454391
rect -46 454351 -34 454385
rect 34 454351 46 454385
rect -46 454345 46 454351
rect -46 454277 46 454283
rect -46 454243 -34 454277
rect 34 454243 46 454277
rect -46 454237 46 454243
rect -102 454193 -56 454205
rect -102 453217 -96 454193
rect -62 453217 -56 454193
rect -102 453205 -56 453217
rect 56 454193 102 454205
rect 56 453217 62 454193
rect 96 453217 102 454193
rect 56 453205 102 453217
rect -46 453167 46 453173
rect -46 453133 -34 453167
rect 34 453133 46 453167
rect -46 453127 46 453133
rect -46 453059 46 453065
rect -46 453025 -34 453059
rect 34 453025 46 453059
rect -46 453019 46 453025
rect -102 452975 -56 452987
rect -102 451999 -96 452975
rect -62 451999 -56 452975
rect -102 451987 -56 451999
rect 56 452975 102 452987
rect 56 451999 62 452975
rect 96 451999 102 452975
rect 56 451987 102 451999
rect -46 451949 46 451955
rect -46 451915 -34 451949
rect 34 451915 46 451949
rect -46 451909 46 451915
rect -46 451841 46 451847
rect -46 451807 -34 451841
rect 34 451807 46 451841
rect -46 451801 46 451807
rect -102 451757 -56 451769
rect -102 450781 -96 451757
rect -62 450781 -56 451757
rect -102 450769 -56 450781
rect 56 451757 102 451769
rect 56 450781 62 451757
rect 96 450781 102 451757
rect 56 450769 102 450781
rect -46 450731 46 450737
rect -46 450697 -34 450731
rect 34 450697 46 450731
rect -46 450691 46 450697
rect -46 450623 46 450629
rect -46 450589 -34 450623
rect 34 450589 46 450623
rect -46 450583 46 450589
rect -102 450539 -56 450551
rect -102 449563 -96 450539
rect -62 449563 -56 450539
rect -102 449551 -56 449563
rect 56 450539 102 450551
rect 56 449563 62 450539
rect 96 449563 102 450539
rect 56 449551 102 449563
rect -46 449513 46 449519
rect -46 449479 -34 449513
rect 34 449479 46 449513
rect -46 449473 46 449479
rect -46 449405 46 449411
rect -46 449371 -34 449405
rect 34 449371 46 449405
rect -46 449365 46 449371
rect -102 449321 -56 449333
rect -102 448345 -96 449321
rect -62 448345 -56 449321
rect -102 448333 -56 448345
rect 56 449321 102 449333
rect 56 448345 62 449321
rect 96 448345 102 449321
rect 56 448333 102 448345
rect -46 448295 46 448301
rect -46 448261 -34 448295
rect 34 448261 46 448295
rect -46 448255 46 448261
rect -46 448187 46 448193
rect -46 448153 -34 448187
rect 34 448153 46 448187
rect -46 448147 46 448153
rect -102 448103 -56 448115
rect -102 447127 -96 448103
rect -62 447127 -56 448103
rect -102 447115 -56 447127
rect 56 448103 102 448115
rect 56 447127 62 448103
rect 96 447127 102 448103
rect 56 447115 102 447127
rect -46 447077 46 447083
rect -46 447043 -34 447077
rect 34 447043 46 447077
rect -46 447037 46 447043
rect -46 446969 46 446975
rect -46 446935 -34 446969
rect 34 446935 46 446969
rect -46 446929 46 446935
rect -102 446885 -56 446897
rect -102 445909 -96 446885
rect -62 445909 -56 446885
rect -102 445897 -56 445909
rect 56 446885 102 446897
rect 56 445909 62 446885
rect 96 445909 102 446885
rect 56 445897 102 445909
rect -46 445859 46 445865
rect -46 445825 -34 445859
rect 34 445825 46 445859
rect -46 445819 46 445825
rect -46 445751 46 445757
rect -46 445717 -34 445751
rect 34 445717 46 445751
rect -46 445711 46 445717
rect -102 445667 -56 445679
rect -102 444691 -96 445667
rect -62 444691 -56 445667
rect -102 444679 -56 444691
rect 56 445667 102 445679
rect 56 444691 62 445667
rect 96 444691 102 445667
rect 56 444679 102 444691
rect -46 444641 46 444647
rect -46 444607 -34 444641
rect 34 444607 46 444641
rect -46 444601 46 444607
rect -46 444533 46 444539
rect -46 444499 -34 444533
rect 34 444499 46 444533
rect -46 444493 46 444499
rect -102 444449 -56 444461
rect -102 443473 -96 444449
rect -62 443473 -56 444449
rect -102 443461 -56 443473
rect 56 444449 102 444461
rect 56 443473 62 444449
rect 96 443473 102 444449
rect 56 443461 102 443473
rect -46 443423 46 443429
rect -46 443389 -34 443423
rect 34 443389 46 443423
rect -46 443383 46 443389
rect -46 443315 46 443321
rect -46 443281 -34 443315
rect 34 443281 46 443315
rect -46 443275 46 443281
rect -102 443231 -56 443243
rect -102 442255 -96 443231
rect -62 442255 -56 443231
rect -102 442243 -56 442255
rect 56 443231 102 443243
rect 56 442255 62 443231
rect 96 442255 102 443231
rect 56 442243 102 442255
rect -46 442205 46 442211
rect -46 442171 -34 442205
rect 34 442171 46 442205
rect -46 442165 46 442171
rect -46 442097 46 442103
rect -46 442063 -34 442097
rect 34 442063 46 442097
rect -46 442057 46 442063
rect -102 442013 -56 442025
rect -102 441037 -96 442013
rect -62 441037 -56 442013
rect -102 441025 -56 441037
rect 56 442013 102 442025
rect 56 441037 62 442013
rect 96 441037 102 442013
rect 56 441025 102 441037
rect -46 440987 46 440993
rect -46 440953 -34 440987
rect 34 440953 46 440987
rect -46 440947 46 440953
rect -46 440879 46 440885
rect -46 440845 -34 440879
rect 34 440845 46 440879
rect -46 440839 46 440845
rect -102 440795 -56 440807
rect -102 439819 -96 440795
rect -62 439819 -56 440795
rect -102 439807 -56 439819
rect 56 440795 102 440807
rect 56 439819 62 440795
rect 96 439819 102 440795
rect 56 439807 102 439819
rect -46 439769 46 439775
rect -46 439735 -34 439769
rect 34 439735 46 439769
rect -46 439729 46 439735
rect -46 439661 46 439667
rect -46 439627 -34 439661
rect 34 439627 46 439661
rect -46 439621 46 439627
rect -102 439577 -56 439589
rect -102 438601 -96 439577
rect -62 438601 -56 439577
rect -102 438589 -56 438601
rect 56 439577 102 439589
rect 56 438601 62 439577
rect 96 438601 102 439577
rect 56 438589 102 438601
rect -46 438551 46 438557
rect -46 438517 -34 438551
rect 34 438517 46 438551
rect -46 438511 46 438517
rect -46 438443 46 438449
rect -46 438409 -34 438443
rect 34 438409 46 438443
rect -46 438403 46 438409
rect -102 438359 -56 438371
rect -102 437383 -96 438359
rect -62 437383 -56 438359
rect -102 437371 -56 437383
rect 56 438359 102 438371
rect 56 437383 62 438359
rect 96 437383 102 438359
rect 56 437371 102 437383
rect -46 437333 46 437339
rect -46 437299 -34 437333
rect 34 437299 46 437333
rect -46 437293 46 437299
rect -46 437225 46 437231
rect -46 437191 -34 437225
rect 34 437191 46 437225
rect -46 437185 46 437191
rect -102 437141 -56 437153
rect -102 436165 -96 437141
rect -62 436165 -56 437141
rect -102 436153 -56 436165
rect 56 437141 102 437153
rect 56 436165 62 437141
rect 96 436165 102 437141
rect 56 436153 102 436165
rect -46 436115 46 436121
rect -46 436081 -34 436115
rect 34 436081 46 436115
rect -46 436075 46 436081
rect -46 436007 46 436013
rect -46 435973 -34 436007
rect 34 435973 46 436007
rect -46 435967 46 435973
rect -102 435923 -56 435935
rect -102 434947 -96 435923
rect -62 434947 -56 435923
rect -102 434935 -56 434947
rect 56 435923 102 435935
rect 56 434947 62 435923
rect 96 434947 102 435923
rect 56 434935 102 434947
rect -46 434897 46 434903
rect -46 434863 -34 434897
rect 34 434863 46 434897
rect -46 434857 46 434863
rect -46 434789 46 434795
rect -46 434755 -34 434789
rect 34 434755 46 434789
rect -46 434749 46 434755
rect -102 434705 -56 434717
rect -102 433729 -96 434705
rect -62 433729 -56 434705
rect -102 433717 -56 433729
rect 56 434705 102 434717
rect 56 433729 62 434705
rect 96 433729 102 434705
rect 56 433717 102 433729
rect -46 433679 46 433685
rect -46 433645 -34 433679
rect 34 433645 46 433679
rect -46 433639 46 433645
rect -46 433571 46 433577
rect -46 433537 -34 433571
rect 34 433537 46 433571
rect -46 433531 46 433537
rect -102 433487 -56 433499
rect -102 432511 -96 433487
rect -62 432511 -56 433487
rect -102 432499 -56 432511
rect 56 433487 102 433499
rect 56 432511 62 433487
rect 96 432511 102 433487
rect 56 432499 102 432511
rect -46 432461 46 432467
rect -46 432427 -34 432461
rect 34 432427 46 432461
rect -46 432421 46 432427
rect -46 432353 46 432359
rect -46 432319 -34 432353
rect 34 432319 46 432353
rect -46 432313 46 432319
rect -102 432269 -56 432281
rect -102 431293 -96 432269
rect -62 431293 -56 432269
rect -102 431281 -56 431293
rect 56 432269 102 432281
rect 56 431293 62 432269
rect 96 431293 102 432269
rect 56 431281 102 431293
rect -46 431243 46 431249
rect -46 431209 -34 431243
rect 34 431209 46 431243
rect -46 431203 46 431209
rect -46 431135 46 431141
rect -46 431101 -34 431135
rect 34 431101 46 431135
rect -46 431095 46 431101
rect -102 431051 -56 431063
rect -102 430075 -96 431051
rect -62 430075 -56 431051
rect -102 430063 -56 430075
rect 56 431051 102 431063
rect 56 430075 62 431051
rect 96 430075 102 431051
rect 56 430063 102 430075
rect -46 430025 46 430031
rect -46 429991 -34 430025
rect 34 429991 46 430025
rect -46 429985 46 429991
rect -46 429917 46 429923
rect -46 429883 -34 429917
rect 34 429883 46 429917
rect -46 429877 46 429883
rect -102 429833 -56 429845
rect -102 428857 -96 429833
rect -62 428857 -56 429833
rect -102 428845 -56 428857
rect 56 429833 102 429845
rect 56 428857 62 429833
rect 96 428857 102 429833
rect 56 428845 102 428857
rect -46 428807 46 428813
rect -46 428773 -34 428807
rect 34 428773 46 428807
rect -46 428767 46 428773
rect -46 428699 46 428705
rect -46 428665 -34 428699
rect 34 428665 46 428699
rect -46 428659 46 428665
rect -102 428615 -56 428627
rect -102 427639 -96 428615
rect -62 427639 -56 428615
rect -102 427627 -56 427639
rect 56 428615 102 428627
rect 56 427639 62 428615
rect 96 427639 102 428615
rect 56 427627 102 427639
rect -46 427589 46 427595
rect -46 427555 -34 427589
rect 34 427555 46 427589
rect -46 427549 46 427555
rect -46 427481 46 427487
rect -46 427447 -34 427481
rect 34 427447 46 427481
rect -46 427441 46 427447
rect -102 427397 -56 427409
rect -102 426421 -96 427397
rect -62 426421 -56 427397
rect -102 426409 -56 426421
rect 56 427397 102 427409
rect 56 426421 62 427397
rect 96 426421 102 427397
rect 56 426409 102 426421
rect -46 426371 46 426377
rect -46 426337 -34 426371
rect 34 426337 46 426371
rect -46 426331 46 426337
rect -46 426263 46 426269
rect -46 426229 -34 426263
rect 34 426229 46 426263
rect -46 426223 46 426229
rect -102 426179 -56 426191
rect -102 425203 -96 426179
rect -62 425203 -56 426179
rect -102 425191 -56 425203
rect 56 426179 102 426191
rect 56 425203 62 426179
rect 96 425203 102 426179
rect 56 425191 102 425203
rect -46 425153 46 425159
rect -46 425119 -34 425153
rect 34 425119 46 425153
rect -46 425113 46 425119
rect -46 425045 46 425051
rect -46 425011 -34 425045
rect 34 425011 46 425045
rect -46 425005 46 425011
rect -102 424961 -56 424973
rect -102 423985 -96 424961
rect -62 423985 -56 424961
rect -102 423973 -56 423985
rect 56 424961 102 424973
rect 56 423985 62 424961
rect 96 423985 102 424961
rect 56 423973 102 423985
rect -46 423935 46 423941
rect -46 423901 -34 423935
rect 34 423901 46 423935
rect -46 423895 46 423901
rect -46 423827 46 423833
rect -46 423793 -34 423827
rect 34 423793 46 423827
rect -46 423787 46 423793
rect -102 423743 -56 423755
rect -102 422767 -96 423743
rect -62 422767 -56 423743
rect -102 422755 -56 422767
rect 56 423743 102 423755
rect 56 422767 62 423743
rect 96 422767 102 423743
rect 56 422755 102 422767
rect -46 422717 46 422723
rect -46 422683 -34 422717
rect 34 422683 46 422717
rect -46 422677 46 422683
rect -46 422609 46 422615
rect -46 422575 -34 422609
rect 34 422575 46 422609
rect -46 422569 46 422575
rect -102 422525 -56 422537
rect -102 421549 -96 422525
rect -62 421549 -56 422525
rect -102 421537 -56 421549
rect 56 422525 102 422537
rect 56 421549 62 422525
rect 96 421549 102 422525
rect 56 421537 102 421549
rect -46 421499 46 421505
rect -46 421465 -34 421499
rect 34 421465 46 421499
rect -46 421459 46 421465
rect -46 421391 46 421397
rect -46 421357 -34 421391
rect 34 421357 46 421391
rect -46 421351 46 421357
rect -102 421307 -56 421319
rect -102 420331 -96 421307
rect -62 420331 -56 421307
rect -102 420319 -56 420331
rect 56 421307 102 421319
rect 56 420331 62 421307
rect 96 420331 102 421307
rect 56 420319 102 420331
rect -46 420281 46 420287
rect -46 420247 -34 420281
rect 34 420247 46 420281
rect -46 420241 46 420247
rect -46 420173 46 420179
rect -46 420139 -34 420173
rect 34 420139 46 420173
rect -46 420133 46 420139
rect -102 420089 -56 420101
rect -102 419113 -96 420089
rect -62 419113 -56 420089
rect -102 419101 -56 419113
rect 56 420089 102 420101
rect 56 419113 62 420089
rect 96 419113 102 420089
rect 56 419101 102 419113
rect -46 419063 46 419069
rect -46 419029 -34 419063
rect 34 419029 46 419063
rect -46 419023 46 419029
rect -46 418955 46 418961
rect -46 418921 -34 418955
rect 34 418921 46 418955
rect -46 418915 46 418921
rect -102 418871 -56 418883
rect -102 417895 -96 418871
rect -62 417895 -56 418871
rect -102 417883 -56 417895
rect 56 418871 102 418883
rect 56 417895 62 418871
rect 96 417895 102 418871
rect 56 417883 102 417895
rect -46 417845 46 417851
rect -46 417811 -34 417845
rect 34 417811 46 417845
rect -46 417805 46 417811
rect -46 417737 46 417743
rect -46 417703 -34 417737
rect 34 417703 46 417737
rect -46 417697 46 417703
rect -102 417653 -56 417665
rect -102 416677 -96 417653
rect -62 416677 -56 417653
rect -102 416665 -56 416677
rect 56 417653 102 417665
rect 56 416677 62 417653
rect 96 416677 102 417653
rect 56 416665 102 416677
rect -46 416627 46 416633
rect -46 416593 -34 416627
rect 34 416593 46 416627
rect -46 416587 46 416593
rect -46 416519 46 416525
rect -46 416485 -34 416519
rect 34 416485 46 416519
rect -46 416479 46 416485
rect -102 416435 -56 416447
rect -102 415459 -96 416435
rect -62 415459 -56 416435
rect -102 415447 -56 415459
rect 56 416435 102 416447
rect 56 415459 62 416435
rect 96 415459 102 416435
rect 56 415447 102 415459
rect -46 415409 46 415415
rect -46 415375 -34 415409
rect 34 415375 46 415409
rect -46 415369 46 415375
rect -46 415301 46 415307
rect -46 415267 -34 415301
rect 34 415267 46 415301
rect -46 415261 46 415267
rect -102 415217 -56 415229
rect -102 414241 -96 415217
rect -62 414241 -56 415217
rect -102 414229 -56 414241
rect 56 415217 102 415229
rect 56 414241 62 415217
rect 96 414241 102 415217
rect 56 414229 102 414241
rect -46 414191 46 414197
rect -46 414157 -34 414191
rect 34 414157 46 414191
rect -46 414151 46 414157
rect -46 414083 46 414089
rect -46 414049 -34 414083
rect 34 414049 46 414083
rect -46 414043 46 414049
rect -102 413999 -56 414011
rect -102 413023 -96 413999
rect -62 413023 -56 413999
rect -102 413011 -56 413023
rect 56 413999 102 414011
rect 56 413023 62 413999
rect 96 413023 102 413999
rect 56 413011 102 413023
rect -46 412973 46 412979
rect -46 412939 -34 412973
rect 34 412939 46 412973
rect -46 412933 46 412939
rect -46 412865 46 412871
rect -46 412831 -34 412865
rect 34 412831 46 412865
rect -46 412825 46 412831
rect -102 412781 -56 412793
rect -102 411805 -96 412781
rect -62 411805 -56 412781
rect -102 411793 -56 411805
rect 56 412781 102 412793
rect 56 411805 62 412781
rect 96 411805 102 412781
rect 56 411793 102 411805
rect -46 411755 46 411761
rect -46 411721 -34 411755
rect 34 411721 46 411755
rect -46 411715 46 411721
rect -46 411647 46 411653
rect -46 411613 -34 411647
rect 34 411613 46 411647
rect -46 411607 46 411613
rect -102 411563 -56 411575
rect -102 410587 -96 411563
rect -62 410587 -56 411563
rect -102 410575 -56 410587
rect 56 411563 102 411575
rect 56 410587 62 411563
rect 96 410587 102 411563
rect 56 410575 102 410587
rect -46 410537 46 410543
rect -46 410503 -34 410537
rect 34 410503 46 410537
rect -46 410497 46 410503
rect -46 410429 46 410435
rect -46 410395 -34 410429
rect 34 410395 46 410429
rect -46 410389 46 410395
rect -102 410345 -56 410357
rect -102 409369 -96 410345
rect -62 409369 -56 410345
rect -102 409357 -56 409369
rect 56 410345 102 410357
rect 56 409369 62 410345
rect 96 409369 102 410345
rect 56 409357 102 409369
rect -46 409319 46 409325
rect -46 409285 -34 409319
rect 34 409285 46 409319
rect -46 409279 46 409285
rect -46 409211 46 409217
rect -46 409177 -34 409211
rect 34 409177 46 409211
rect -46 409171 46 409177
rect -102 409127 -56 409139
rect -102 408151 -96 409127
rect -62 408151 -56 409127
rect -102 408139 -56 408151
rect 56 409127 102 409139
rect 56 408151 62 409127
rect 96 408151 102 409127
rect 56 408139 102 408151
rect -46 408101 46 408107
rect -46 408067 -34 408101
rect 34 408067 46 408101
rect -46 408061 46 408067
rect -46 407993 46 407999
rect -46 407959 -34 407993
rect 34 407959 46 407993
rect -46 407953 46 407959
rect -102 407909 -56 407921
rect -102 406933 -96 407909
rect -62 406933 -56 407909
rect -102 406921 -56 406933
rect 56 407909 102 407921
rect 56 406933 62 407909
rect 96 406933 102 407909
rect 56 406921 102 406933
rect -46 406883 46 406889
rect -46 406849 -34 406883
rect 34 406849 46 406883
rect -46 406843 46 406849
rect -46 406775 46 406781
rect -46 406741 -34 406775
rect 34 406741 46 406775
rect -46 406735 46 406741
rect -102 406691 -56 406703
rect -102 405715 -96 406691
rect -62 405715 -56 406691
rect -102 405703 -56 405715
rect 56 406691 102 406703
rect 56 405715 62 406691
rect 96 405715 102 406691
rect 56 405703 102 405715
rect -46 405665 46 405671
rect -46 405631 -34 405665
rect 34 405631 46 405665
rect -46 405625 46 405631
rect -46 405557 46 405563
rect -46 405523 -34 405557
rect 34 405523 46 405557
rect -46 405517 46 405523
rect -102 405473 -56 405485
rect -102 404497 -96 405473
rect -62 404497 -56 405473
rect -102 404485 -56 404497
rect 56 405473 102 405485
rect 56 404497 62 405473
rect 96 404497 102 405473
rect 56 404485 102 404497
rect -46 404447 46 404453
rect -46 404413 -34 404447
rect 34 404413 46 404447
rect -46 404407 46 404413
rect -46 404339 46 404345
rect -46 404305 -34 404339
rect 34 404305 46 404339
rect -46 404299 46 404305
rect -102 404255 -56 404267
rect -102 403279 -96 404255
rect -62 403279 -56 404255
rect -102 403267 -56 403279
rect 56 404255 102 404267
rect 56 403279 62 404255
rect 96 403279 102 404255
rect 56 403267 102 403279
rect -46 403229 46 403235
rect -46 403195 -34 403229
rect 34 403195 46 403229
rect -46 403189 46 403195
rect -46 403121 46 403127
rect -46 403087 -34 403121
rect 34 403087 46 403121
rect -46 403081 46 403087
rect -102 403037 -56 403049
rect -102 402061 -96 403037
rect -62 402061 -56 403037
rect -102 402049 -56 402061
rect 56 403037 102 403049
rect 56 402061 62 403037
rect 96 402061 102 403037
rect 56 402049 102 402061
rect -46 402011 46 402017
rect -46 401977 -34 402011
rect 34 401977 46 402011
rect -46 401971 46 401977
rect -46 401903 46 401909
rect -46 401869 -34 401903
rect 34 401869 46 401903
rect -46 401863 46 401869
rect -102 401819 -56 401831
rect -102 400843 -96 401819
rect -62 400843 -56 401819
rect -102 400831 -56 400843
rect 56 401819 102 401831
rect 56 400843 62 401819
rect 96 400843 102 401819
rect 56 400831 102 400843
rect -46 400793 46 400799
rect -46 400759 -34 400793
rect 34 400759 46 400793
rect -46 400753 46 400759
rect -46 400685 46 400691
rect -46 400651 -34 400685
rect 34 400651 46 400685
rect -46 400645 46 400651
rect -102 400601 -56 400613
rect -102 399625 -96 400601
rect -62 399625 -56 400601
rect -102 399613 -56 399625
rect 56 400601 102 400613
rect 56 399625 62 400601
rect 96 399625 102 400601
rect 56 399613 102 399625
rect -46 399575 46 399581
rect -46 399541 -34 399575
rect 34 399541 46 399575
rect -46 399535 46 399541
rect -46 399467 46 399473
rect -46 399433 -34 399467
rect 34 399433 46 399467
rect -46 399427 46 399433
rect -102 399383 -56 399395
rect -102 398407 -96 399383
rect -62 398407 -56 399383
rect -102 398395 -56 398407
rect 56 399383 102 399395
rect 56 398407 62 399383
rect 96 398407 102 399383
rect 56 398395 102 398407
rect -46 398357 46 398363
rect -46 398323 -34 398357
rect 34 398323 46 398357
rect -46 398317 46 398323
rect -46 398249 46 398255
rect -46 398215 -34 398249
rect 34 398215 46 398249
rect -46 398209 46 398215
rect -102 398165 -56 398177
rect -102 397189 -96 398165
rect -62 397189 -56 398165
rect -102 397177 -56 397189
rect 56 398165 102 398177
rect 56 397189 62 398165
rect 96 397189 102 398165
rect 56 397177 102 397189
rect -46 397139 46 397145
rect -46 397105 -34 397139
rect 34 397105 46 397139
rect -46 397099 46 397105
rect -46 397031 46 397037
rect -46 396997 -34 397031
rect 34 396997 46 397031
rect -46 396991 46 396997
rect -102 396947 -56 396959
rect -102 395971 -96 396947
rect -62 395971 -56 396947
rect -102 395959 -56 395971
rect 56 396947 102 396959
rect 56 395971 62 396947
rect 96 395971 102 396947
rect 56 395959 102 395971
rect -46 395921 46 395927
rect -46 395887 -34 395921
rect 34 395887 46 395921
rect -46 395881 46 395887
rect -46 395813 46 395819
rect -46 395779 -34 395813
rect 34 395779 46 395813
rect -46 395773 46 395779
rect -102 395729 -56 395741
rect -102 394753 -96 395729
rect -62 394753 -56 395729
rect -102 394741 -56 394753
rect 56 395729 102 395741
rect 56 394753 62 395729
rect 96 394753 102 395729
rect 56 394741 102 394753
rect -46 394703 46 394709
rect -46 394669 -34 394703
rect 34 394669 46 394703
rect -46 394663 46 394669
rect -46 394595 46 394601
rect -46 394561 -34 394595
rect 34 394561 46 394595
rect -46 394555 46 394561
rect -102 394511 -56 394523
rect -102 393535 -96 394511
rect -62 393535 -56 394511
rect -102 393523 -56 393535
rect 56 394511 102 394523
rect 56 393535 62 394511
rect 96 393535 102 394511
rect 56 393523 102 393535
rect -46 393485 46 393491
rect -46 393451 -34 393485
rect 34 393451 46 393485
rect -46 393445 46 393451
rect -46 393377 46 393383
rect -46 393343 -34 393377
rect 34 393343 46 393377
rect -46 393337 46 393343
rect -102 393293 -56 393305
rect -102 392317 -96 393293
rect -62 392317 -56 393293
rect -102 392305 -56 392317
rect 56 393293 102 393305
rect 56 392317 62 393293
rect 96 392317 102 393293
rect 56 392305 102 392317
rect -46 392267 46 392273
rect -46 392233 -34 392267
rect 34 392233 46 392267
rect -46 392227 46 392233
rect -46 392159 46 392165
rect -46 392125 -34 392159
rect 34 392125 46 392159
rect -46 392119 46 392125
rect -102 392075 -56 392087
rect -102 391099 -96 392075
rect -62 391099 -56 392075
rect -102 391087 -56 391099
rect 56 392075 102 392087
rect 56 391099 62 392075
rect 96 391099 102 392075
rect 56 391087 102 391099
rect -46 391049 46 391055
rect -46 391015 -34 391049
rect 34 391015 46 391049
rect -46 391009 46 391015
rect -46 390941 46 390947
rect -46 390907 -34 390941
rect 34 390907 46 390941
rect -46 390901 46 390907
rect -102 390857 -56 390869
rect -102 389881 -96 390857
rect -62 389881 -56 390857
rect -102 389869 -56 389881
rect 56 390857 102 390869
rect 56 389881 62 390857
rect 96 389881 102 390857
rect 56 389869 102 389881
rect -46 389831 46 389837
rect -46 389797 -34 389831
rect 34 389797 46 389831
rect -46 389791 46 389797
rect -46 389723 46 389729
rect -46 389689 -34 389723
rect 34 389689 46 389723
rect -46 389683 46 389689
rect -102 389639 -56 389651
rect -102 388663 -96 389639
rect -62 388663 -56 389639
rect -102 388651 -56 388663
rect 56 389639 102 389651
rect 56 388663 62 389639
rect 96 388663 102 389639
rect 56 388651 102 388663
rect -46 388613 46 388619
rect -46 388579 -34 388613
rect 34 388579 46 388613
rect -46 388573 46 388579
rect -46 388505 46 388511
rect -46 388471 -34 388505
rect 34 388471 46 388505
rect -46 388465 46 388471
rect -102 388421 -56 388433
rect -102 387445 -96 388421
rect -62 387445 -56 388421
rect -102 387433 -56 387445
rect 56 388421 102 388433
rect 56 387445 62 388421
rect 96 387445 102 388421
rect 56 387433 102 387445
rect -46 387395 46 387401
rect -46 387361 -34 387395
rect 34 387361 46 387395
rect -46 387355 46 387361
rect -46 387287 46 387293
rect -46 387253 -34 387287
rect 34 387253 46 387287
rect -46 387247 46 387253
rect -102 387203 -56 387215
rect -102 386227 -96 387203
rect -62 386227 -56 387203
rect -102 386215 -56 386227
rect 56 387203 102 387215
rect 56 386227 62 387203
rect 96 386227 102 387203
rect 56 386215 102 386227
rect -46 386177 46 386183
rect -46 386143 -34 386177
rect 34 386143 46 386177
rect -46 386137 46 386143
rect -46 386069 46 386075
rect -46 386035 -34 386069
rect 34 386035 46 386069
rect -46 386029 46 386035
rect -102 385985 -56 385997
rect -102 385009 -96 385985
rect -62 385009 -56 385985
rect -102 384997 -56 385009
rect 56 385985 102 385997
rect 56 385009 62 385985
rect 96 385009 102 385985
rect 56 384997 102 385009
rect -46 384959 46 384965
rect -46 384925 -34 384959
rect 34 384925 46 384959
rect -46 384919 46 384925
rect -46 384851 46 384857
rect -46 384817 -34 384851
rect 34 384817 46 384851
rect -46 384811 46 384817
rect -102 384767 -56 384779
rect -102 383791 -96 384767
rect -62 383791 -56 384767
rect -102 383779 -56 383791
rect 56 384767 102 384779
rect 56 383791 62 384767
rect 96 383791 102 384767
rect 56 383779 102 383791
rect -46 383741 46 383747
rect -46 383707 -34 383741
rect 34 383707 46 383741
rect -46 383701 46 383707
rect -46 383633 46 383639
rect -46 383599 -34 383633
rect 34 383599 46 383633
rect -46 383593 46 383599
rect -102 383549 -56 383561
rect -102 382573 -96 383549
rect -62 382573 -56 383549
rect -102 382561 -56 382573
rect 56 383549 102 383561
rect 56 382573 62 383549
rect 96 382573 102 383549
rect 56 382561 102 382573
rect -46 382523 46 382529
rect -46 382489 -34 382523
rect 34 382489 46 382523
rect -46 382483 46 382489
rect -46 382415 46 382421
rect -46 382381 -34 382415
rect 34 382381 46 382415
rect -46 382375 46 382381
rect -102 382331 -56 382343
rect -102 381355 -96 382331
rect -62 381355 -56 382331
rect -102 381343 -56 381355
rect 56 382331 102 382343
rect 56 381355 62 382331
rect 96 381355 102 382331
rect 56 381343 102 381355
rect -46 381305 46 381311
rect -46 381271 -34 381305
rect 34 381271 46 381305
rect -46 381265 46 381271
rect -46 381197 46 381203
rect -46 381163 -34 381197
rect 34 381163 46 381197
rect -46 381157 46 381163
rect -102 381113 -56 381125
rect -102 380137 -96 381113
rect -62 380137 -56 381113
rect -102 380125 -56 380137
rect 56 381113 102 381125
rect 56 380137 62 381113
rect 96 380137 102 381113
rect 56 380125 102 380137
rect -46 380087 46 380093
rect -46 380053 -34 380087
rect 34 380053 46 380087
rect -46 380047 46 380053
rect -46 379979 46 379985
rect -46 379945 -34 379979
rect 34 379945 46 379979
rect -46 379939 46 379945
rect -102 379895 -56 379907
rect -102 378919 -96 379895
rect -62 378919 -56 379895
rect -102 378907 -56 378919
rect 56 379895 102 379907
rect 56 378919 62 379895
rect 96 378919 102 379895
rect 56 378907 102 378919
rect -46 378869 46 378875
rect -46 378835 -34 378869
rect 34 378835 46 378869
rect -46 378829 46 378835
rect -46 378761 46 378767
rect -46 378727 -34 378761
rect 34 378727 46 378761
rect -46 378721 46 378727
rect -102 378677 -56 378689
rect -102 377701 -96 378677
rect -62 377701 -56 378677
rect -102 377689 -56 377701
rect 56 378677 102 378689
rect 56 377701 62 378677
rect 96 377701 102 378677
rect 56 377689 102 377701
rect -46 377651 46 377657
rect -46 377617 -34 377651
rect 34 377617 46 377651
rect -46 377611 46 377617
rect -46 377543 46 377549
rect -46 377509 -34 377543
rect 34 377509 46 377543
rect -46 377503 46 377509
rect -102 377459 -56 377471
rect -102 376483 -96 377459
rect -62 376483 -56 377459
rect -102 376471 -56 376483
rect 56 377459 102 377471
rect 56 376483 62 377459
rect 96 376483 102 377459
rect 56 376471 102 376483
rect -46 376433 46 376439
rect -46 376399 -34 376433
rect 34 376399 46 376433
rect -46 376393 46 376399
rect -46 376325 46 376331
rect -46 376291 -34 376325
rect 34 376291 46 376325
rect -46 376285 46 376291
rect -102 376241 -56 376253
rect -102 375265 -96 376241
rect -62 375265 -56 376241
rect -102 375253 -56 375265
rect 56 376241 102 376253
rect 56 375265 62 376241
rect 96 375265 102 376241
rect 56 375253 102 375265
rect -46 375215 46 375221
rect -46 375181 -34 375215
rect 34 375181 46 375215
rect -46 375175 46 375181
rect -46 375107 46 375113
rect -46 375073 -34 375107
rect 34 375073 46 375107
rect -46 375067 46 375073
rect -102 375023 -56 375035
rect -102 374047 -96 375023
rect -62 374047 -56 375023
rect -102 374035 -56 374047
rect 56 375023 102 375035
rect 56 374047 62 375023
rect 96 374047 102 375023
rect 56 374035 102 374047
rect -46 373997 46 374003
rect -46 373963 -34 373997
rect 34 373963 46 373997
rect -46 373957 46 373963
rect -46 373889 46 373895
rect -46 373855 -34 373889
rect 34 373855 46 373889
rect -46 373849 46 373855
rect -102 373805 -56 373817
rect -102 372829 -96 373805
rect -62 372829 -56 373805
rect -102 372817 -56 372829
rect 56 373805 102 373817
rect 56 372829 62 373805
rect 96 372829 102 373805
rect 56 372817 102 372829
rect -46 372779 46 372785
rect -46 372745 -34 372779
rect 34 372745 46 372779
rect -46 372739 46 372745
rect -46 372671 46 372677
rect -46 372637 -34 372671
rect 34 372637 46 372671
rect -46 372631 46 372637
rect -102 372587 -56 372599
rect -102 371611 -96 372587
rect -62 371611 -56 372587
rect -102 371599 -56 371611
rect 56 372587 102 372599
rect 56 371611 62 372587
rect 96 371611 102 372587
rect 56 371599 102 371611
rect -46 371561 46 371567
rect -46 371527 -34 371561
rect 34 371527 46 371561
rect -46 371521 46 371527
rect -46 371453 46 371459
rect -46 371419 -34 371453
rect 34 371419 46 371453
rect -46 371413 46 371419
rect -102 371369 -56 371381
rect -102 370393 -96 371369
rect -62 370393 -56 371369
rect -102 370381 -56 370393
rect 56 371369 102 371381
rect 56 370393 62 371369
rect 96 370393 102 371369
rect 56 370381 102 370393
rect -46 370343 46 370349
rect -46 370309 -34 370343
rect 34 370309 46 370343
rect -46 370303 46 370309
rect -46 370235 46 370241
rect -46 370201 -34 370235
rect 34 370201 46 370235
rect -46 370195 46 370201
rect -102 370151 -56 370163
rect -102 369175 -96 370151
rect -62 369175 -56 370151
rect -102 369163 -56 369175
rect 56 370151 102 370163
rect 56 369175 62 370151
rect 96 369175 102 370151
rect 56 369163 102 369175
rect -46 369125 46 369131
rect -46 369091 -34 369125
rect 34 369091 46 369125
rect -46 369085 46 369091
rect -46 369017 46 369023
rect -46 368983 -34 369017
rect 34 368983 46 369017
rect -46 368977 46 368983
rect -102 368933 -56 368945
rect -102 367957 -96 368933
rect -62 367957 -56 368933
rect -102 367945 -56 367957
rect 56 368933 102 368945
rect 56 367957 62 368933
rect 96 367957 102 368933
rect 56 367945 102 367957
rect -46 367907 46 367913
rect -46 367873 -34 367907
rect 34 367873 46 367907
rect -46 367867 46 367873
rect -46 367799 46 367805
rect -46 367765 -34 367799
rect 34 367765 46 367799
rect -46 367759 46 367765
rect -102 367715 -56 367727
rect -102 366739 -96 367715
rect -62 366739 -56 367715
rect -102 366727 -56 366739
rect 56 367715 102 367727
rect 56 366739 62 367715
rect 96 366739 102 367715
rect 56 366727 102 366739
rect -46 366689 46 366695
rect -46 366655 -34 366689
rect 34 366655 46 366689
rect -46 366649 46 366655
rect -46 366581 46 366587
rect -46 366547 -34 366581
rect 34 366547 46 366581
rect -46 366541 46 366547
rect -102 366497 -56 366509
rect -102 365521 -96 366497
rect -62 365521 -56 366497
rect -102 365509 -56 365521
rect 56 366497 102 366509
rect 56 365521 62 366497
rect 96 365521 102 366497
rect 56 365509 102 365521
rect -46 365471 46 365477
rect -46 365437 -34 365471
rect 34 365437 46 365471
rect -46 365431 46 365437
rect -46 365363 46 365369
rect -46 365329 -34 365363
rect 34 365329 46 365363
rect -46 365323 46 365329
rect -102 365279 -56 365291
rect -102 364303 -96 365279
rect -62 364303 -56 365279
rect -102 364291 -56 364303
rect 56 365279 102 365291
rect 56 364303 62 365279
rect 96 364303 102 365279
rect 56 364291 102 364303
rect -46 364253 46 364259
rect -46 364219 -34 364253
rect 34 364219 46 364253
rect -46 364213 46 364219
rect -46 364145 46 364151
rect -46 364111 -34 364145
rect 34 364111 46 364145
rect -46 364105 46 364111
rect -102 364061 -56 364073
rect -102 363085 -96 364061
rect -62 363085 -56 364061
rect -102 363073 -56 363085
rect 56 364061 102 364073
rect 56 363085 62 364061
rect 96 363085 102 364061
rect 56 363073 102 363085
rect -46 363035 46 363041
rect -46 363001 -34 363035
rect 34 363001 46 363035
rect -46 362995 46 363001
rect -46 362927 46 362933
rect -46 362893 -34 362927
rect 34 362893 46 362927
rect -46 362887 46 362893
rect -102 362843 -56 362855
rect -102 361867 -96 362843
rect -62 361867 -56 362843
rect -102 361855 -56 361867
rect 56 362843 102 362855
rect 56 361867 62 362843
rect 96 361867 102 362843
rect 56 361855 102 361867
rect -46 361817 46 361823
rect -46 361783 -34 361817
rect 34 361783 46 361817
rect -46 361777 46 361783
rect -46 361709 46 361715
rect -46 361675 -34 361709
rect 34 361675 46 361709
rect -46 361669 46 361675
rect -102 361625 -56 361637
rect -102 360649 -96 361625
rect -62 360649 -56 361625
rect -102 360637 -56 360649
rect 56 361625 102 361637
rect 56 360649 62 361625
rect 96 360649 102 361625
rect 56 360637 102 360649
rect -46 360599 46 360605
rect -46 360565 -34 360599
rect 34 360565 46 360599
rect -46 360559 46 360565
rect -46 360491 46 360497
rect -46 360457 -34 360491
rect 34 360457 46 360491
rect -46 360451 46 360457
rect -102 360407 -56 360419
rect -102 359431 -96 360407
rect -62 359431 -56 360407
rect -102 359419 -56 359431
rect 56 360407 102 360419
rect 56 359431 62 360407
rect 96 359431 102 360407
rect 56 359419 102 359431
rect -46 359381 46 359387
rect -46 359347 -34 359381
rect 34 359347 46 359381
rect -46 359341 46 359347
rect -46 359273 46 359279
rect -46 359239 -34 359273
rect 34 359239 46 359273
rect -46 359233 46 359239
rect -102 359189 -56 359201
rect -102 358213 -96 359189
rect -62 358213 -56 359189
rect -102 358201 -56 358213
rect 56 359189 102 359201
rect 56 358213 62 359189
rect 96 358213 102 359189
rect 56 358201 102 358213
rect -46 358163 46 358169
rect -46 358129 -34 358163
rect 34 358129 46 358163
rect -46 358123 46 358129
rect -46 358055 46 358061
rect -46 358021 -34 358055
rect 34 358021 46 358055
rect -46 358015 46 358021
rect -102 357971 -56 357983
rect -102 356995 -96 357971
rect -62 356995 -56 357971
rect -102 356983 -56 356995
rect 56 357971 102 357983
rect 56 356995 62 357971
rect 96 356995 102 357971
rect 56 356983 102 356995
rect -46 356945 46 356951
rect -46 356911 -34 356945
rect 34 356911 46 356945
rect -46 356905 46 356911
rect -46 356837 46 356843
rect -46 356803 -34 356837
rect 34 356803 46 356837
rect -46 356797 46 356803
rect -102 356753 -56 356765
rect -102 355777 -96 356753
rect -62 355777 -56 356753
rect -102 355765 -56 355777
rect 56 356753 102 356765
rect 56 355777 62 356753
rect 96 355777 102 356753
rect 56 355765 102 355777
rect -46 355727 46 355733
rect -46 355693 -34 355727
rect 34 355693 46 355727
rect -46 355687 46 355693
rect -46 355619 46 355625
rect -46 355585 -34 355619
rect 34 355585 46 355619
rect -46 355579 46 355585
rect -102 355535 -56 355547
rect -102 354559 -96 355535
rect -62 354559 -56 355535
rect -102 354547 -56 354559
rect 56 355535 102 355547
rect 56 354559 62 355535
rect 96 354559 102 355535
rect 56 354547 102 354559
rect -46 354509 46 354515
rect -46 354475 -34 354509
rect 34 354475 46 354509
rect -46 354469 46 354475
rect -46 354401 46 354407
rect -46 354367 -34 354401
rect 34 354367 46 354401
rect -46 354361 46 354367
rect -102 354317 -56 354329
rect -102 353341 -96 354317
rect -62 353341 -56 354317
rect -102 353329 -56 353341
rect 56 354317 102 354329
rect 56 353341 62 354317
rect 96 353341 102 354317
rect 56 353329 102 353341
rect -46 353291 46 353297
rect -46 353257 -34 353291
rect 34 353257 46 353291
rect -46 353251 46 353257
rect -46 353183 46 353189
rect -46 353149 -34 353183
rect 34 353149 46 353183
rect -46 353143 46 353149
rect -102 353099 -56 353111
rect -102 352123 -96 353099
rect -62 352123 -56 353099
rect -102 352111 -56 352123
rect 56 353099 102 353111
rect 56 352123 62 353099
rect 96 352123 102 353099
rect 56 352111 102 352123
rect -46 352073 46 352079
rect -46 352039 -34 352073
rect 34 352039 46 352073
rect -46 352033 46 352039
rect -46 351965 46 351971
rect -46 351931 -34 351965
rect 34 351931 46 351965
rect -46 351925 46 351931
rect -102 351881 -56 351893
rect -102 350905 -96 351881
rect -62 350905 -56 351881
rect -102 350893 -56 350905
rect 56 351881 102 351893
rect 56 350905 62 351881
rect 96 350905 102 351881
rect 56 350893 102 350905
rect -46 350855 46 350861
rect -46 350821 -34 350855
rect 34 350821 46 350855
rect -46 350815 46 350821
rect -46 350747 46 350753
rect -46 350713 -34 350747
rect 34 350713 46 350747
rect -46 350707 46 350713
rect -102 350663 -56 350675
rect -102 349687 -96 350663
rect -62 349687 -56 350663
rect -102 349675 -56 349687
rect 56 350663 102 350675
rect 56 349687 62 350663
rect 96 349687 102 350663
rect 56 349675 102 349687
rect -46 349637 46 349643
rect -46 349603 -34 349637
rect 34 349603 46 349637
rect -46 349597 46 349603
rect -46 349529 46 349535
rect -46 349495 -34 349529
rect 34 349495 46 349529
rect -46 349489 46 349495
rect -102 349445 -56 349457
rect -102 348469 -96 349445
rect -62 348469 -56 349445
rect -102 348457 -56 348469
rect 56 349445 102 349457
rect 56 348469 62 349445
rect 96 348469 102 349445
rect 56 348457 102 348469
rect -46 348419 46 348425
rect -46 348385 -34 348419
rect 34 348385 46 348419
rect -46 348379 46 348385
rect -46 348311 46 348317
rect -46 348277 -34 348311
rect 34 348277 46 348311
rect -46 348271 46 348277
rect -102 348227 -56 348239
rect -102 347251 -96 348227
rect -62 347251 -56 348227
rect -102 347239 -56 347251
rect 56 348227 102 348239
rect 56 347251 62 348227
rect 96 347251 102 348227
rect 56 347239 102 347251
rect -46 347201 46 347207
rect -46 347167 -34 347201
rect 34 347167 46 347201
rect -46 347161 46 347167
rect -46 347093 46 347099
rect -46 347059 -34 347093
rect 34 347059 46 347093
rect -46 347053 46 347059
rect -102 347009 -56 347021
rect -102 346033 -96 347009
rect -62 346033 -56 347009
rect -102 346021 -56 346033
rect 56 347009 102 347021
rect 56 346033 62 347009
rect 96 346033 102 347009
rect 56 346021 102 346033
rect -46 345983 46 345989
rect -46 345949 -34 345983
rect 34 345949 46 345983
rect -46 345943 46 345949
rect -46 345875 46 345881
rect -46 345841 -34 345875
rect 34 345841 46 345875
rect -46 345835 46 345841
rect -102 345791 -56 345803
rect -102 344815 -96 345791
rect -62 344815 -56 345791
rect -102 344803 -56 344815
rect 56 345791 102 345803
rect 56 344815 62 345791
rect 96 344815 102 345791
rect 56 344803 102 344815
rect -46 344765 46 344771
rect -46 344731 -34 344765
rect 34 344731 46 344765
rect -46 344725 46 344731
rect -46 344657 46 344663
rect -46 344623 -34 344657
rect 34 344623 46 344657
rect -46 344617 46 344623
rect -102 344573 -56 344585
rect -102 343597 -96 344573
rect -62 343597 -56 344573
rect -102 343585 -56 343597
rect 56 344573 102 344585
rect 56 343597 62 344573
rect 96 343597 102 344573
rect 56 343585 102 343597
rect -46 343547 46 343553
rect -46 343513 -34 343547
rect 34 343513 46 343547
rect -46 343507 46 343513
rect -46 343439 46 343445
rect -46 343405 -34 343439
rect 34 343405 46 343439
rect -46 343399 46 343405
rect -102 343355 -56 343367
rect -102 342379 -96 343355
rect -62 342379 -56 343355
rect -102 342367 -56 342379
rect 56 343355 102 343367
rect 56 342379 62 343355
rect 96 342379 102 343355
rect 56 342367 102 342379
rect -46 342329 46 342335
rect -46 342295 -34 342329
rect 34 342295 46 342329
rect -46 342289 46 342295
rect -46 342221 46 342227
rect -46 342187 -34 342221
rect 34 342187 46 342221
rect -46 342181 46 342187
rect -102 342137 -56 342149
rect -102 341161 -96 342137
rect -62 341161 -56 342137
rect -102 341149 -56 341161
rect 56 342137 102 342149
rect 56 341161 62 342137
rect 96 341161 102 342137
rect 56 341149 102 341161
rect -46 341111 46 341117
rect -46 341077 -34 341111
rect 34 341077 46 341111
rect -46 341071 46 341077
rect -46 341003 46 341009
rect -46 340969 -34 341003
rect 34 340969 46 341003
rect -46 340963 46 340969
rect -102 340919 -56 340931
rect -102 339943 -96 340919
rect -62 339943 -56 340919
rect -102 339931 -56 339943
rect 56 340919 102 340931
rect 56 339943 62 340919
rect 96 339943 102 340919
rect 56 339931 102 339943
rect -46 339893 46 339899
rect -46 339859 -34 339893
rect 34 339859 46 339893
rect -46 339853 46 339859
rect -46 339785 46 339791
rect -46 339751 -34 339785
rect 34 339751 46 339785
rect -46 339745 46 339751
rect -102 339701 -56 339713
rect -102 338725 -96 339701
rect -62 338725 -56 339701
rect -102 338713 -56 338725
rect 56 339701 102 339713
rect 56 338725 62 339701
rect 96 338725 102 339701
rect 56 338713 102 338725
rect -46 338675 46 338681
rect -46 338641 -34 338675
rect 34 338641 46 338675
rect -46 338635 46 338641
rect -46 338567 46 338573
rect -46 338533 -34 338567
rect 34 338533 46 338567
rect -46 338527 46 338533
rect -102 338483 -56 338495
rect -102 337507 -96 338483
rect -62 337507 -56 338483
rect -102 337495 -56 337507
rect 56 338483 102 338495
rect 56 337507 62 338483
rect 96 337507 102 338483
rect 56 337495 102 337507
rect -46 337457 46 337463
rect -46 337423 -34 337457
rect 34 337423 46 337457
rect -46 337417 46 337423
rect -46 337349 46 337355
rect -46 337315 -34 337349
rect 34 337315 46 337349
rect -46 337309 46 337315
rect -102 337265 -56 337277
rect -102 336289 -96 337265
rect -62 336289 -56 337265
rect -102 336277 -56 336289
rect 56 337265 102 337277
rect 56 336289 62 337265
rect 96 336289 102 337265
rect 56 336277 102 336289
rect -46 336239 46 336245
rect -46 336205 -34 336239
rect 34 336205 46 336239
rect -46 336199 46 336205
rect -46 336131 46 336137
rect -46 336097 -34 336131
rect 34 336097 46 336131
rect -46 336091 46 336097
rect -102 336047 -56 336059
rect -102 335071 -96 336047
rect -62 335071 -56 336047
rect -102 335059 -56 335071
rect 56 336047 102 336059
rect 56 335071 62 336047
rect 96 335071 102 336047
rect 56 335059 102 335071
rect -46 335021 46 335027
rect -46 334987 -34 335021
rect 34 334987 46 335021
rect -46 334981 46 334987
rect -46 334913 46 334919
rect -46 334879 -34 334913
rect 34 334879 46 334913
rect -46 334873 46 334879
rect -102 334829 -56 334841
rect -102 333853 -96 334829
rect -62 333853 -56 334829
rect -102 333841 -56 333853
rect 56 334829 102 334841
rect 56 333853 62 334829
rect 96 333853 102 334829
rect 56 333841 102 333853
rect -46 333803 46 333809
rect -46 333769 -34 333803
rect 34 333769 46 333803
rect -46 333763 46 333769
rect -46 333695 46 333701
rect -46 333661 -34 333695
rect 34 333661 46 333695
rect -46 333655 46 333661
rect -102 333611 -56 333623
rect -102 332635 -96 333611
rect -62 332635 -56 333611
rect -102 332623 -56 332635
rect 56 333611 102 333623
rect 56 332635 62 333611
rect 96 332635 102 333611
rect 56 332623 102 332635
rect -46 332585 46 332591
rect -46 332551 -34 332585
rect 34 332551 46 332585
rect -46 332545 46 332551
rect -46 332477 46 332483
rect -46 332443 -34 332477
rect 34 332443 46 332477
rect -46 332437 46 332443
rect -102 332393 -56 332405
rect -102 331417 -96 332393
rect -62 331417 -56 332393
rect -102 331405 -56 331417
rect 56 332393 102 332405
rect 56 331417 62 332393
rect 96 331417 102 332393
rect 56 331405 102 331417
rect -46 331367 46 331373
rect -46 331333 -34 331367
rect 34 331333 46 331367
rect -46 331327 46 331333
rect -46 331259 46 331265
rect -46 331225 -34 331259
rect 34 331225 46 331259
rect -46 331219 46 331225
rect -102 331175 -56 331187
rect -102 330199 -96 331175
rect -62 330199 -56 331175
rect -102 330187 -56 330199
rect 56 331175 102 331187
rect 56 330199 62 331175
rect 96 330199 102 331175
rect 56 330187 102 330199
rect -46 330149 46 330155
rect -46 330115 -34 330149
rect 34 330115 46 330149
rect -46 330109 46 330115
rect -46 330041 46 330047
rect -46 330007 -34 330041
rect 34 330007 46 330041
rect -46 330001 46 330007
rect -102 329957 -56 329969
rect -102 328981 -96 329957
rect -62 328981 -56 329957
rect -102 328969 -56 328981
rect 56 329957 102 329969
rect 56 328981 62 329957
rect 96 328981 102 329957
rect 56 328969 102 328981
rect -46 328931 46 328937
rect -46 328897 -34 328931
rect 34 328897 46 328931
rect -46 328891 46 328897
rect -46 328823 46 328829
rect -46 328789 -34 328823
rect 34 328789 46 328823
rect -46 328783 46 328789
rect -102 328739 -56 328751
rect -102 327763 -96 328739
rect -62 327763 -56 328739
rect -102 327751 -56 327763
rect 56 328739 102 328751
rect 56 327763 62 328739
rect 96 327763 102 328739
rect 56 327751 102 327763
rect -46 327713 46 327719
rect -46 327679 -34 327713
rect 34 327679 46 327713
rect -46 327673 46 327679
rect -46 327605 46 327611
rect -46 327571 -34 327605
rect 34 327571 46 327605
rect -46 327565 46 327571
rect -102 327521 -56 327533
rect -102 326545 -96 327521
rect -62 326545 -56 327521
rect -102 326533 -56 326545
rect 56 327521 102 327533
rect 56 326545 62 327521
rect 96 326545 102 327521
rect 56 326533 102 326545
rect -46 326495 46 326501
rect -46 326461 -34 326495
rect 34 326461 46 326495
rect -46 326455 46 326461
rect -46 326387 46 326393
rect -46 326353 -34 326387
rect 34 326353 46 326387
rect -46 326347 46 326353
rect -102 326303 -56 326315
rect -102 325327 -96 326303
rect -62 325327 -56 326303
rect -102 325315 -56 325327
rect 56 326303 102 326315
rect 56 325327 62 326303
rect 96 325327 102 326303
rect 56 325315 102 325327
rect -46 325277 46 325283
rect -46 325243 -34 325277
rect 34 325243 46 325277
rect -46 325237 46 325243
rect -46 325169 46 325175
rect -46 325135 -34 325169
rect 34 325135 46 325169
rect -46 325129 46 325135
rect -102 325085 -56 325097
rect -102 324109 -96 325085
rect -62 324109 -56 325085
rect -102 324097 -56 324109
rect 56 325085 102 325097
rect 56 324109 62 325085
rect 96 324109 102 325085
rect 56 324097 102 324109
rect -46 324059 46 324065
rect -46 324025 -34 324059
rect 34 324025 46 324059
rect -46 324019 46 324025
rect -46 323951 46 323957
rect -46 323917 -34 323951
rect 34 323917 46 323951
rect -46 323911 46 323917
rect -102 323867 -56 323879
rect -102 322891 -96 323867
rect -62 322891 -56 323867
rect -102 322879 -56 322891
rect 56 323867 102 323879
rect 56 322891 62 323867
rect 96 322891 102 323867
rect 56 322879 102 322891
rect -46 322841 46 322847
rect -46 322807 -34 322841
rect 34 322807 46 322841
rect -46 322801 46 322807
rect -46 322733 46 322739
rect -46 322699 -34 322733
rect 34 322699 46 322733
rect -46 322693 46 322699
rect -102 322649 -56 322661
rect -102 321673 -96 322649
rect -62 321673 -56 322649
rect -102 321661 -56 321673
rect 56 322649 102 322661
rect 56 321673 62 322649
rect 96 321673 102 322649
rect 56 321661 102 321673
rect -46 321623 46 321629
rect -46 321589 -34 321623
rect 34 321589 46 321623
rect -46 321583 46 321589
rect -46 321515 46 321521
rect -46 321481 -34 321515
rect 34 321481 46 321515
rect -46 321475 46 321481
rect -102 321431 -56 321443
rect -102 320455 -96 321431
rect -62 320455 -56 321431
rect -102 320443 -56 320455
rect 56 321431 102 321443
rect 56 320455 62 321431
rect 96 320455 102 321431
rect 56 320443 102 320455
rect -46 320405 46 320411
rect -46 320371 -34 320405
rect 34 320371 46 320405
rect -46 320365 46 320371
rect -46 320297 46 320303
rect -46 320263 -34 320297
rect 34 320263 46 320297
rect -46 320257 46 320263
rect -102 320213 -56 320225
rect -102 319237 -96 320213
rect -62 319237 -56 320213
rect -102 319225 -56 319237
rect 56 320213 102 320225
rect 56 319237 62 320213
rect 96 319237 102 320213
rect 56 319225 102 319237
rect -46 319187 46 319193
rect -46 319153 -34 319187
rect 34 319153 46 319187
rect -46 319147 46 319153
rect -46 319079 46 319085
rect -46 319045 -34 319079
rect 34 319045 46 319079
rect -46 319039 46 319045
rect -102 318995 -56 319007
rect -102 318019 -96 318995
rect -62 318019 -56 318995
rect -102 318007 -56 318019
rect 56 318995 102 319007
rect 56 318019 62 318995
rect 96 318019 102 318995
rect 56 318007 102 318019
rect -46 317969 46 317975
rect -46 317935 -34 317969
rect 34 317935 46 317969
rect -46 317929 46 317935
rect -46 317861 46 317867
rect -46 317827 -34 317861
rect 34 317827 46 317861
rect -46 317821 46 317827
rect -102 317777 -56 317789
rect -102 316801 -96 317777
rect -62 316801 -56 317777
rect -102 316789 -56 316801
rect 56 317777 102 317789
rect 56 316801 62 317777
rect 96 316801 102 317777
rect 56 316789 102 316801
rect -46 316751 46 316757
rect -46 316717 -34 316751
rect 34 316717 46 316751
rect -46 316711 46 316717
rect -46 316643 46 316649
rect -46 316609 -34 316643
rect 34 316609 46 316643
rect -46 316603 46 316609
rect -102 316559 -56 316571
rect -102 315583 -96 316559
rect -62 315583 -56 316559
rect -102 315571 -56 315583
rect 56 316559 102 316571
rect 56 315583 62 316559
rect 96 315583 102 316559
rect 56 315571 102 315583
rect -46 315533 46 315539
rect -46 315499 -34 315533
rect 34 315499 46 315533
rect -46 315493 46 315499
rect -46 315425 46 315431
rect -46 315391 -34 315425
rect 34 315391 46 315425
rect -46 315385 46 315391
rect -102 315341 -56 315353
rect -102 314365 -96 315341
rect -62 314365 -56 315341
rect -102 314353 -56 314365
rect 56 315341 102 315353
rect 56 314365 62 315341
rect 96 314365 102 315341
rect 56 314353 102 314365
rect -46 314315 46 314321
rect -46 314281 -34 314315
rect 34 314281 46 314315
rect -46 314275 46 314281
rect -46 314207 46 314213
rect -46 314173 -34 314207
rect 34 314173 46 314207
rect -46 314167 46 314173
rect -102 314123 -56 314135
rect -102 313147 -96 314123
rect -62 313147 -56 314123
rect -102 313135 -56 313147
rect 56 314123 102 314135
rect 56 313147 62 314123
rect 96 313147 102 314123
rect 56 313135 102 313147
rect -46 313097 46 313103
rect -46 313063 -34 313097
rect 34 313063 46 313097
rect -46 313057 46 313063
rect -46 312989 46 312995
rect -46 312955 -34 312989
rect 34 312955 46 312989
rect -46 312949 46 312955
rect -102 312905 -56 312917
rect -102 311929 -96 312905
rect -62 311929 -56 312905
rect -102 311917 -56 311929
rect 56 312905 102 312917
rect 56 311929 62 312905
rect 96 311929 102 312905
rect 56 311917 102 311929
rect -46 311879 46 311885
rect -46 311845 -34 311879
rect 34 311845 46 311879
rect -46 311839 46 311845
rect -46 311771 46 311777
rect -46 311737 -34 311771
rect 34 311737 46 311771
rect -46 311731 46 311737
rect -102 311687 -56 311699
rect -102 310711 -96 311687
rect -62 310711 -56 311687
rect -102 310699 -56 310711
rect 56 311687 102 311699
rect 56 310711 62 311687
rect 96 310711 102 311687
rect 56 310699 102 310711
rect -46 310661 46 310667
rect -46 310627 -34 310661
rect 34 310627 46 310661
rect -46 310621 46 310627
rect -46 310553 46 310559
rect -46 310519 -34 310553
rect 34 310519 46 310553
rect -46 310513 46 310519
rect -102 310469 -56 310481
rect -102 309493 -96 310469
rect -62 309493 -56 310469
rect -102 309481 -56 309493
rect 56 310469 102 310481
rect 56 309493 62 310469
rect 96 309493 102 310469
rect 56 309481 102 309493
rect -46 309443 46 309449
rect -46 309409 -34 309443
rect 34 309409 46 309443
rect -46 309403 46 309409
rect -46 309335 46 309341
rect -46 309301 -34 309335
rect 34 309301 46 309335
rect -46 309295 46 309301
rect -102 309251 -56 309263
rect -102 308275 -96 309251
rect -62 308275 -56 309251
rect -102 308263 -56 308275
rect 56 309251 102 309263
rect 56 308275 62 309251
rect 96 308275 102 309251
rect 56 308263 102 308275
rect -46 308225 46 308231
rect -46 308191 -34 308225
rect 34 308191 46 308225
rect -46 308185 46 308191
rect -46 308117 46 308123
rect -46 308083 -34 308117
rect 34 308083 46 308117
rect -46 308077 46 308083
rect -102 308033 -56 308045
rect -102 307057 -96 308033
rect -62 307057 -56 308033
rect -102 307045 -56 307057
rect 56 308033 102 308045
rect 56 307057 62 308033
rect 96 307057 102 308033
rect 56 307045 102 307057
rect -46 307007 46 307013
rect -46 306973 -34 307007
rect 34 306973 46 307007
rect -46 306967 46 306973
rect -46 306899 46 306905
rect -46 306865 -34 306899
rect 34 306865 46 306899
rect -46 306859 46 306865
rect -102 306815 -56 306827
rect -102 305839 -96 306815
rect -62 305839 -56 306815
rect -102 305827 -56 305839
rect 56 306815 102 306827
rect 56 305839 62 306815
rect 96 305839 102 306815
rect 56 305827 102 305839
rect -46 305789 46 305795
rect -46 305755 -34 305789
rect 34 305755 46 305789
rect -46 305749 46 305755
rect -46 305681 46 305687
rect -46 305647 -34 305681
rect 34 305647 46 305681
rect -46 305641 46 305647
rect -102 305597 -56 305609
rect -102 304621 -96 305597
rect -62 304621 -56 305597
rect -102 304609 -56 304621
rect 56 305597 102 305609
rect 56 304621 62 305597
rect 96 304621 102 305597
rect 56 304609 102 304621
rect -46 304571 46 304577
rect -46 304537 -34 304571
rect 34 304537 46 304571
rect -46 304531 46 304537
rect -46 304463 46 304469
rect -46 304429 -34 304463
rect 34 304429 46 304463
rect -46 304423 46 304429
rect -102 304379 -56 304391
rect -102 303403 -96 304379
rect -62 303403 -56 304379
rect -102 303391 -56 303403
rect 56 304379 102 304391
rect 56 303403 62 304379
rect 96 303403 102 304379
rect 56 303391 102 303403
rect -46 303353 46 303359
rect -46 303319 -34 303353
rect 34 303319 46 303353
rect -46 303313 46 303319
rect -46 303245 46 303251
rect -46 303211 -34 303245
rect 34 303211 46 303245
rect -46 303205 46 303211
rect -102 303161 -56 303173
rect -102 302185 -96 303161
rect -62 302185 -56 303161
rect -102 302173 -56 302185
rect 56 303161 102 303173
rect 56 302185 62 303161
rect 96 302185 102 303161
rect 56 302173 102 302185
rect -46 302135 46 302141
rect -46 302101 -34 302135
rect 34 302101 46 302135
rect -46 302095 46 302101
rect -46 302027 46 302033
rect -46 301993 -34 302027
rect 34 301993 46 302027
rect -46 301987 46 301993
rect -102 301943 -56 301955
rect -102 300967 -96 301943
rect -62 300967 -56 301943
rect -102 300955 -56 300967
rect 56 301943 102 301955
rect 56 300967 62 301943
rect 96 300967 102 301943
rect 56 300955 102 300967
rect -46 300917 46 300923
rect -46 300883 -34 300917
rect 34 300883 46 300917
rect -46 300877 46 300883
rect -46 300809 46 300815
rect -46 300775 -34 300809
rect 34 300775 46 300809
rect -46 300769 46 300775
rect -102 300725 -56 300737
rect -102 299749 -96 300725
rect -62 299749 -56 300725
rect -102 299737 -56 299749
rect 56 300725 102 300737
rect 56 299749 62 300725
rect 96 299749 102 300725
rect 56 299737 102 299749
rect -46 299699 46 299705
rect -46 299665 -34 299699
rect 34 299665 46 299699
rect -46 299659 46 299665
rect -46 299591 46 299597
rect -46 299557 -34 299591
rect 34 299557 46 299591
rect -46 299551 46 299557
rect -102 299507 -56 299519
rect -102 298531 -96 299507
rect -62 298531 -56 299507
rect -102 298519 -56 298531
rect 56 299507 102 299519
rect 56 298531 62 299507
rect 96 298531 102 299507
rect 56 298519 102 298531
rect -46 298481 46 298487
rect -46 298447 -34 298481
rect 34 298447 46 298481
rect -46 298441 46 298447
rect -46 298373 46 298379
rect -46 298339 -34 298373
rect 34 298339 46 298373
rect -46 298333 46 298339
rect -102 298289 -56 298301
rect -102 297313 -96 298289
rect -62 297313 -56 298289
rect -102 297301 -56 297313
rect 56 298289 102 298301
rect 56 297313 62 298289
rect 96 297313 102 298289
rect 56 297301 102 297313
rect -46 297263 46 297269
rect -46 297229 -34 297263
rect 34 297229 46 297263
rect -46 297223 46 297229
rect -46 297155 46 297161
rect -46 297121 -34 297155
rect 34 297121 46 297155
rect -46 297115 46 297121
rect -102 297071 -56 297083
rect -102 296095 -96 297071
rect -62 296095 -56 297071
rect -102 296083 -56 296095
rect 56 297071 102 297083
rect 56 296095 62 297071
rect 96 296095 102 297071
rect 56 296083 102 296095
rect -46 296045 46 296051
rect -46 296011 -34 296045
rect 34 296011 46 296045
rect -46 296005 46 296011
rect -46 295937 46 295943
rect -46 295903 -34 295937
rect 34 295903 46 295937
rect -46 295897 46 295903
rect -102 295853 -56 295865
rect -102 294877 -96 295853
rect -62 294877 -56 295853
rect -102 294865 -56 294877
rect 56 295853 102 295865
rect 56 294877 62 295853
rect 96 294877 102 295853
rect 56 294865 102 294877
rect -46 294827 46 294833
rect -46 294793 -34 294827
rect 34 294793 46 294827
rect -46 294787 46 294793
rect -46 294719 46 294725
rect -46 294685 -34 294719
rect 34 294685 46 294719
rect -46 294679 46 294685
rect -102 294635 -56 294647
rect -102 293659 -96 294635
rect -62 293659 -56 294635
rect -102 293647 -56 293659
rect 56 294635 102 294647
rect 56 293659 62 294635
rect 96 293659 102 294635
rect 56 293647 102 293659
rect -46 293609 46 293615
rect -46 293575 -34 293609
rect 34 293575 46 293609
rect -46 293569 46 293575
rect -46 293501 46 293507
rect -46 293467 -34 293501
rect 34 293467 46 293501
rect -46 293461 46 293467
rect -102 293417 -56 293429
rect -102 292441 -96 293417
rect -62 292441 -56 293417
rect -102 292429 -56 292441
rect 56 293417 102 293429
rect 56 292441 62 293417
rect 96 292441 102 293417
rect 56 292429 102 292441
rect -46 292391 46 292397
rect -46 292357 -34 292391
rect 34 292357 46 292391
rect -46 292351 46 292357
rect -46 292283 46 292289
rect -46 292249 -34 292283
rect 34 292249 46 292283
rect -46 292243 46 292249
rect -102 292199 -56 292211
rect -102 291223 -96 292199
rect -62 291223 -56 292199
rect -102 291211 -56 291223
rect 56 292199 102 292211
rect 56 291223 62 292199
rect 96 291223 102 292199
rect 56 291211 102 291223
rect -46 291173 46 291179
rect -46 291139 -34 291173
rect 34 291139 46 291173
rect -46 291133 46 291139
rect -46 291065 46 291071
rect -46 291031 -34 291065
rect 34 291031 46 291065
rect -46 291025 46 291031
rect -102 290981 -56 290993
rect -102 290005 -96 290981
rect -62 290005 -56 290981
rect -102 289993 -56 290005
rect 56 290981 102 290993
rect 56 290005 62 290981
rect 96 290005 102 290981
rect 56 289993 102 290005
rect -46 289955 46 289961
rect -46 289921 -34 289955
rect 34 289921 46 289955
rect -46 289915 46 289921
rect -46 289847 46 289853
rect -46 289813 -34 289847
rect 34 289813 46 289847
rect -46 289807 46 289813
rect -102 289763 -56 289775
rect -102 288787 -96 289763
rect -62 288787 -56 289763
rect -102 288775 -56 288787
rect 56 289763 102 289775
rect 56 288787 62 289763
rect 96 288787 102 289763
rect 56 288775 102 288787
rect -46 288737 46 288743
rect -46 288703 -34 288737
rect 34 288703 46 288737
rect -46 288697 46 288703
rect -46 288629 46 288635
rect -46 288595 -34 288629
rect 34 288595 46 288629
rect -46 288589 46 288595
rect -102 288545 -56 288557
rect -102 287569 -96 288545
rect -62 287569 -56 288545
rect -102 287557 -56 287569
rect 56 288545 102 288557
rect 56 287569 62 288545
rect 96 287569 102 288545
rect 56 287557 102 287569
rect -46 287519 46 287525
rect -46 287485 -34 287519
rect 34 287485 46 287519
rect -46 287479 46 287485
rect -46 287411 46 287417
rect -46 287377 -34 287411
rect 34 287377 46 287411
rect -46 287371 46 287377
rect -102 287327 -56 287339
rect -102 286351 -96 287327
rect -62 286351 -56 287327
rect -102 286339 -56 286351
rect 56 287327 102 287339
rect 56 286351 62 287327
rect 96 286351 102 287327
rect 56 286339 102 286351
rect -46 286301 46 286307
rect -46 286267 -34 286301
rect 34 286267 46 286301
rect -46 286261 46 286267
rect -46 286193 46 286199
rect -46 286159 -34 286193
rect 34 286159 46 286193
rect -46 286153 46 286159
rect -102 286109 -56 286121
rect -102 285133 -96 286109
rect -62 285133 -56 286109
rect -102 285121 -56 285133
rect 56 286109 102 286121
rect 56 285133 62 286109
rect 96 285133 102 286109
rect 56 285121 102 285133
rect -46 285083 46 285089
rect -46 285049 -34 285083
rect 34 285049 46 285083
rect -46 285043 46 285049
rect -46 284975 46 284981
rect -46 284941 -34 284975
rect 34 284941 46 284975
rect -46 284935 46 284941
rect -102 284891 -56 284903
rect -102 283915 -96 284891
rect -62 283915 -56 284891
rect -102 283903 -56 283915
rect 56 284891 102 284903
rect 56 283915 62 284891
rect 96 283915 102 284891
rect 56 283903 102 283915
rect -46 283865 46 283871
rect -46 283831 -34 283865
rect 34 283831 46 283865
rect -46 283825 46 283831
rect -46 283757 46 283763
rect -46 283723 -34 283757
rect 34 283723 46 283757
rect -46 283717 46 283723
rect -102 283673 -56 283685
rect -102 282697 -96 283673
rect -62 282697 -56 283673
rect -102 282685 -56 282697
rect 56 283673 102 283685
rect 56 282697 62 283673
rect 96 282697 102 283673
rect 56 282685 102 282697
rect -46 282647 46 282653
rect -46 282613 -34 282647
rect 34 282613 46 282647
rect -46 282607 46 282613
rect -46 282539 46 282545
rect -46 282505 -34 282539
rect 34 282505 46 282539
rect -46 282499 46 282505
rect -102 282455 -56 282467
rect -102 281479 -96 282455
rect -62 281479 -56 282455
rect -102 281467 -56 281479
rect 56 282455 102 282467
rect 56 281479 62 282455
rect 96 281479 102 282455
rect 56 281467 102 281479
rect -46 281429 46 281435
rect -46 281395 -34 281429
rect 34 281395 46 281429
rect -46 281389 46 281395
rect -46 281321 46 281327
rect -46 281287 -34 281321
rect 34 281287 46 281321
rect -46 281281 46 281287
rect -102 281237 -56 281249
rect -102 280261 -96 281237
rect -62 280261 -56 281237
rect -102 280249 -56 280261
rect 56 281237 102 281249
rect 56 280261 62 281237
rect 96 280261 102 281237
rect 56 280249 102 280261
rect -46 280211 46 280217
rect -46 280177 -34 280211
rect 34 280177 46 280211
rect -46 280171 46 280177
rect -46 280103 46 280109
rect -46 280069 -34 280103
rect 34 280069 46 280103
rect -46 280063 46 280069
rect -102 280019 -56 280031
rect -102 279043 -96 280019
rect -62 279043 -56 280019
rect -102 279031 -56 279043
rect 56 280019 102 280031
rect 56 279043 62 280019
rect 96 279043 102 280019
rect 56 279031 102 279043
rect -46 278993 46 278999
rect -46 278959 -34 278993
rect 34 278959 46 278993
rect -46 278953 46 278959
rect -46 278885 46 278891
rect -46 278851 -34 278885
rect 34 278851 46 278885
rect -46 278845 46 278851
rect -102 278801 -56 278813
rect -102 277825 -96 278801
rect -62 277825 -56 278801
rect -102 277813 -56 277825
rect 56 278801 102 278813
rect 56 277825 62 278801
rect 96 277825 102 278801
rect 56 277813 102 277825
rect -46 277775 46 277781
rect -46 277741 -34 277775
rect 34 277741 46 277775
rect -46 277735 46 277741
rect -46 277667 46 277673
rect -46 277633 -34 277667
rect 34 277633 46 277667
rect -46 277627 46 277633
rect -102 277583 -56 277595
rect -102 276607 -96 277583
rect -62 276607 -56 277583
rect -102 276595 -56 276607
rect 56 277583 102 277595
rect 56 276607 62 277583
rect 96 276607 102 277583
rect 56 276595 102 276607
rect -46 276557 46 276563
rect -46 276523 -34 276557
rect 34 276523 46 276557
rect -46 276517 46 276523
rect -46 276449 46 276455
rect -46 276415 -34 276449
rect 34 276415 46 276449
rect -46 276409 46 276415
rect -102 276365 -56 276377
rect -102 275389 -96 276365
rect -62 275389 -56 276365
rect -102 275377 -56 275389
rect 56 276365 102 276377
rect 56 275389 62 276365
rect 96 275389 102 276365
rect 56 275377 102 275389
rect -46 275339 46 275345
rect -46 275305 -34 275339
rect 34 275305 46 275339
rect -46 275299 46 275305
rect -46 275231 46 275237
rect -46 275197 -34 275231
rect 34 275197 46 275231
rect -46 275191 46 275197
rect -102 275147 -56 275159
rect -102 274171 -96 275147
rect -62 274171 -56 275147
rect -102 274159 -56 274171
rect 56 275147 102 275159
rect 56 274171 62 275147
rect 96 274171 102 275147
rect 56 274159 102 274171
rect -46 274121 46 274127
rect -46 274087 -34 274121
rect 34 274087 46 274121
rect -46 274081 46 274087
rect -46 274013 46 274019
rect -46 273979 -34 274013
rect 34 273979 46 274013
rect -46 273973 46 273979
rect -102 273929 -56 273941
rect -102 272953 -96 273929
rect -62 272953 -56 273929
rect -102 272941 -56 272953
rect 56 273929 102 273941
rect 56 272953 62 273929
rect 96 272953 102 273929
rect 56 272941 102 272953
rect -46 272903 46 272909
rect -46 272869 -34 272903
rect 34 272869 46 272903
rect -46 272863 46 272869
rect -46 272795 46 272801
rect -46 272761 -34 272795
rect 34 272761 46 272795
rect -46 272755 46 272761
rect -102 272711 -56 272723
rect -102 271735 -96 272711
rect -62 271735 -56 272711
rect -102 271723 -56 271735
rect 56 272711 102 272723
rect 56 271735 62 272711
rect 96 271735 102 272711
rect 56 271723 102 271735
rect -46 271685 46 271691
rect -46 271651 -34 271685
rect 34 271651 46 271685
rect -46 271645 46 271651
rect -46 271577 46 271583
rect -46 271543 -34 271577
rect 34 271543 46 271577
rect -46 271537 46 271543
rect -102 271493 -56 271505
rect -102 270517 -96 271493
rect -62 270517 -56 271493
rect -102 270505 -56 270517
rect 56 271493 102 271505
rect 56 270517 62 271493
rect 96 270517 102 271493
rect 56 270505 102 270517
rect -46 270467 46 270473
rect -46 270433 -34 270467
rect 34 270433 46 270467
rect -46 270427 46 270433
rect -46 270359 46 270365
rect -46 270325 -34 270359
rect 34 270325 46 270359
rect -46 270319 46 270325
rect -102 270275 -56 270287
rect -102 269299 -96 270275
rect -62 269299 -56 270275
rect -102 269287 -56 269299
rect 56 270275 102 270287
rect 56 269299 62 270275
rect 96 269299 102 270275
rect 56 269287 102 269299
rect -46 269249 46 269255
rect -46 269215 -34 269249
rect 34 269215 46 269249
rect -46 269209 46 269215
rect -46 269141 46 269147
rect -46 269107 -34 269141
rect 34 269107 46 269141
rect -46 269101 46 269107
rect -102 269057 -56 269069
rect -102 268081 -96 269057
rect -62 268081 -56 269057
rect -102 268069 -56 268081
rect 56 269057 102 269069
rect 56 268081 62 269057
rect 96 268081 102 269057
rect 56 268069 102 268081
rect -46 268031 46 268037
rect -46 267997 -34 268031
rect 34 267997 46 268031
rect -46 267991 46 267997
rect -46 267923 46 267929
rect -46 267889 -34 267923
rect 34 267889 46 267923
rect -46 267883 46 267889
rect -102 267839 -56 267851
rect -102 266863 -96 267839
rect -62 266863 -56 267839
rect -102 266851 -56 266863
rect 56 267839 102 267851
rect 56 266863 62 267839
rect 96 266863 102 267839
rect 56 266851 102 266863
rect -46 266813 46 266819
rect -46 266779 -34 266813
rect 34 266779 46 266813
rect -46 266773 46 266779
rect -46 266705 46 266711
rect -46 266671 -34 266705
rect 34 266671 46 266705
rect -46 266665 46 266671
rect -102 266621 -56 266633
rect -102 265645 -96 266621
rect -62 265645 -56 266621
rect -102 265633 -56 265645
rect 56 266621 102 266633
rect 56 265645 62 266621
rect 96 265645 102 266621
rect 56 265633 102 265645
rect -46 265595 46 265601
rect -46 265561 -34 265595
rect 34 265561 46 265595
rect -46 265555 46 265561
rect -46 265487 46 265493
rect -46 265453 -34 265487
rect 34 265453 46 265487
rect -46 265447 46 265453
rect -102 265403 -56 265415
rect -102 264427 -96 265403
rect -62 264427 -56 265403
rect -102 264415 -56 264427
rect 56 265403 102 265415
rect 56 264427 62 265403
rect 96 264427 102 265403
rect 56 264415 102 264427
rect -46 264377 46 264383
rect -46 264343 -34 264377
rect 34 264343 46 264377
rect -46 264337 46 264343
rect -46 264269 46 264275
rect -46 264235 -34 264269
rect 34 264235 46 264269
rect -46 264229 46 264235
rect -102 264185 -56 264197
rect -102 263209 -96 264185
rect -62 263209 -56 264185
rect -102 263197 -56 263209
rect 56 264185 102 264197
rect 56 263209 62 264185
rect 96 263209 102 264185
rect 56 263197 102 263209
rect -46 263159 46 263165
rect -46 263125 -34 263159
rect 34 263125 46 263159
rect -46 263119 46 263125
rect -46 263051 46 263057
rect -46 263017 -34 263051
rect 34 263017 46 263051
rect -46 263011 46 263017
rect -102 262967 -56 262979
rect -102 261991 -96 262967
rect -62 261991 -56 262967
rect -102 261979 -56 261991
rect 56 262967 102 262979
rect 56 261991 62 262967
rect 96 261991 102 262967
rect 56 261979 102 261991
rect -46 261941 46 261947
rect -46 261907 -34 261941
rect 34 261907 46 261941
rect -46 261901 46 261907
rect -46 261833 46 261839
rect -46 261799 -34 261833
rect 34 261799 46 261833
rect -46 261793 46 261799
rect -102 261749 -56 261761
rect -102 260773 -96 261749
rect -62 260773 -56 261749
rect -102 260761 -56 260773
rect 56 261749 102 261761
rect 56 260773 62 261749
rect 96 260773 102 261749
rect 56 260761 102 260773
rect -46 260723 46 260729
rect -46 260689 -34 260723
rect 34 260689 46 260723
rect -46 260683 46 260689
rect -46 260615 46 260621
rect -46 260581 -34 260615
rect 34 260581 46 260615
rect -46 260575 46 260581
rect -102 260531 -56 260543
rect -102 259555 -96 260531
rect -62 259555 -56 260531
rect -102 259543 -56 259555
rect 56 260531 102 260543
rect 56 259555 62 260531
rect 96 259555 102 260531
rect 56 259543 102 259555
rect -46 259505 46 259511
rect -46 259471 -34 259505
rect 34 259471 46 259505
rect -46 259465 46 259471
rect -46 259397 46 259403
rect -46 259363 -34 259397
rect 34 259363 46 259397
rect -46 259357 46 259363
rect -102 259313 -56 259325
rect -102 258337 -96 259313
rect -62 258337 -56 259313
rect -102 258325 -56 258337
rect 56 259313 102 259325
rect 56 258337 62 259313
rect 96 258337 102 259313
rect 56 258325 102 258337
rect -46 258287 46 258293
rect -46 258253 -34 258287
rect 34 258253 46 258287
rect -46 258247 46 258253
rect -46 258179 46 258185
rect -46 258145 -34 258179
rect 34 258145 46 258179
rect -46 258139 46 258145
rect -102 258095 -56 258107
rect -102 257119 -96 258095
rect -62 257119 -56 258095
rect -102 257107 -56 257119
rect 56 258095 102 258107
rect 56 257119 62 258095
rect 96 257119 102 258095
rect 56 257107 102 257119
rect -46 257069 46 257075
rect -46 257035 -34 257069
rect 34 257035 46 257069
rect -46 257029 46 257035
rect -46 256961 46 256967
rect -46 256927 -34 256961
rect 34 256927 46 256961
rect -46 256921 46 256927
rect -102 256877 -56 256889
rect -102 255901 -96 256877
rect -62 255901 -56 256877
rect -102 255889 -56 255901
rect 56 256877 102 256889
rect 56 255901 62 256877
rect 96 255901 102 256877
rect 56 255889 102 255901
rect -46 255851 46 255857
rect -46 255817 -34 255851
rect 34 255817 46 255851
rect -46 255811 46 255817
rect -46 255743 46 255749
rect -46 255709 -34 255743
rect 34 255709 46 255743
rect -46 255703 46 255709
rect -102 255659 -56 255671
rect -102 254683 -96 255659
rect -62 254683 -56 255659
rect -102 254671 -56 254683
rect 56 255659 102 255671
rect 56 254683 62 255659
rect 96 254683 102 255659
rect 56 254671 102 254683
rect -46 254633 46 254639
rect -46 254599 -34 254633
rect 34 254599 46 254633
rect -46 254593 46 254599
rect -46 254525 46 254531
rect -46 254491 -34 254525
rect 34 254491 46 254525
rect -46 254485 46 254491
rect -102 254441 -56 254453
rect -102 253465 -96 254441
rect -62 253465 -56 254441
rect -102 253453 -56 253465
rect 56 254441 102 254453
rect 56 253465 62 254441
rect 96 253465 102 254441
rect 56 253453 102 253465
rect -46 253415 46 253421
rect -46 253381 -34 253415
rect 34 253381 46 253415
rect -46 253375 46 253381
rect -46 253307 46 253313
rect -46 253273 -34 253307
rect 34 253273 46 253307
rect -46 253267 46 253273
rect -102 253223 -56 253235
rect -102 252247 -96 253223
rect -62 252247 -56 253223
rect -102 252235 -56 252247
rect 56 253223 102 253235
rect 56 252247 62 253223
rect 96 252247 102 253223
rect 56 252235 102 252247
rect -46 252197 46 252203
rect -46 252163 -34 252197
rect 34 252163 46 252197
rect -46 252157 46 252163
rect -46 252089 46 252095
rect -46 252055 -34 252089
rect 34 252055 46 252089
rect -46 252049 46 252055
rect -102 252005 -56 252017
rect -102 251029 -96 252005
rect -62 251029 -56 252005
rect -102 251017 -56 251029
rect 56 252005 102 252017
rect 56 251029 62 252005
rect 96 251029 102 252005
rect 56 251017 102 251029
rect -46 250979 46 250985
rect -46 250945 -34 250979
rect 34 250945 46 250979
rect -46 250939 46 250945
rect -46 250871 46 250877
rect -46 250837 -34 250871
rect 34 250837 46 250871
rect -46 250831 46 250837
rect -102 250787 -56 250799
rect -102 249811 -96 250787
rect -62 249811 -56 250787
rect -102 249799 -56 249811
rect 56 250787 102 250799
rect 56 249811 62 250787
rect 96 249811 102 250787
rect 56 249799 102 249811
rect -46 249761 46 249767
rect -46 249727 -34 249761
rect 34 249727 46 249761
rect -46 249721 46 249727
rect -46 249653 46 249659
rect -46 249619 -34 249653
rect 34 249619 46 249653
rect -46 249613 46 249619
rect -102 249569 -56 249581
rect -102 248593 -96 249569
rect -62 248593 -56 249569
rect -102 248581 -56 248593
rect 56 249569 102 249581
rect 56 248593 62 249569
rect 96 248593 102 249569
rect 56 248581 102 248593
rect -46 248543 46 248549
rect -46 248509 -34 248543
rect 34 248509 46 248543
rect -46 248503 46 248509
rect -46 248435 46 248441
rect -46 248401 -34 248435
rect 34 248401 46 248435
rect -46 248395 46 248401
rect -102 248351 -56 248363
rect -102 247375 -96 248351
rect -62 247375 -56 248351
rect -102 247363 -56 247375
rect 56 248351 102 248363
rect 56 247375 62 248351
rect 96 247375 102 248351
rect 56 247363 102 247375
rect -46 247325 46 247331
rect -46 247291 -34 247325
rect 34 247291 46 247325
rect -46 247285 46 247291
rect -46 247217 46 247223
rect -46 247183 -34 247217
rect 34 247183 46 247217
rect -46 247177 46 247183
rect -102 247133 -56 247145
rect -102 246157 -96 247133
rect -62 246157 -56 247133
rect -102 246145 -56 246157
rect 56 247133 102 247145
rect 56 246157 62 247133
rect 96 246157 102 247133
rect 56 246145 102 246157
rect -46 246107 46 246113
rect -46 246073 -34 246107
rect 34 246073 46 246107
rect -46 246067 46 246073
rect -46 245999 46 246005
rect -46 245965 -34 245999
rect 34 245965 46 245999
rect -46 245959 46 245965
rect -102 245915 -56 245927
rect -102 244939 -96 245915
rect -62 244939 -56 245915
rect -102 244927 -56 244939
rect 56 245915 102 245927
rect 56 244939 62 245915
rect 96 244939 102 245915
rect 56 244927 102 244939
rect -46 244889 46 244895
rect -46 244855 -34 244889
rect 34 244855 46 244889
rect -46 244849 46 244855
rect -46 244781 46 244787
rect -46 244747 -34 244781
rect 34 244747 46 244781
rect -46 244741 46 244747
rect -102 244697 -56 244709
rect -102 243721 -96 244697
rect -62 243721 -56 244697
rect -102 243709 -56 243721
rect 56 244697 102 244709
rect 56 243721 62 244697
rect 96 243721 102 244697
rect 56 243709 102 243721
rect -46 243671 46 243677
rect -46 243637 -34 243671
rect 34 243637 46 243671
rect -46 243631 46 243637
rect -46 243563 46 243569
rect -46 243529 -34 243563
rect 34 243529 46 243563
rect -46 243523 46 243529
rect -102 243479 -56 243491
rect -102 242503 -96 243479
rect -62 242503 -56 243479
rect -102 242491 -56 242503
rect 56 243479 102 243491
rect 56 242503 62 243479
rect 96 242503 102 243479
rect 56 242491 102 242503
rect -46 242453 46 242459
rect -46 242419 -34 242453
rect 34 242419 46 242453
rect -46 242413 46 242419
rect -46 242345 46 242351
rect -46 242311 -34 242345
rect 34 242311 46 242345
rect -46 242305 46 242311
rect -102 242261 -56 242273
rect -102 241285 -96 242261
rect -62 241285 -56 242261
rect -102 241273 -56 241285
rect 56 242261 102 242273
rect 56 241285 62 242261
rect 96 241285 102 242261
rect 56 241273 102 241285
rect -46 241235 46 241241
rect -46 241201 -34 241235
rect 34 241201 46 241235
rect -46 241195 46 241201
rect -46 241127 46 241133
rect -46 241093 -34 241127
rect 34 241093 46 241127
rect -46 241087 46 241093
rect -102 241043 -56 241055
rect -102 240067 -96 241043
rect -62 240067 -56 241043
rect -102 240055 -56 240067
rect 56 241043 102 241055
rect 56 240067 62 241043
rect 96 240067 102 241043
rect 56 240055 102 240067
rect -46 240017 46 240023
rect -46 239983 -34 240017
rect 34 239983 46 240017
rect -46 239977 46 239983
rect -46 239909 46 239915
rect -46 239875 -34 239909
rect 34 239875 46 239909
rect -46 239869 46 239875
rect -102 239825 -56 239837
rect -102 238849 -96 239825
rect -62 238849 -56 239825
rect -102 238837 -56 238849
rect 56 239825 102 239837
rect 56 238849 62 239825
rect 96 238849 102 239825
rect 56 238837 102 238849
rect -46 238799 46 238805
rect -46 238765 -34 238799
rect 34 238765 46 238799
rect -46 238759 46 238765
rect -46 238691 46 238697
rect -46 238657 -34 238691
rect 34 238657 46 238691
rect -46 238651 46 238657
rect -102 238607 -56 238619
rect -102 237631 -96 238607
rect -62 237631 -56 238607
rect -102 237619 -56 237631
rect 56 238607 102 238619
rect 56 237631 62 238607
rect 96 237631 102 238607
rect 56 237619 102 237631
rect -46 237581 46 237587
rect -46 237547 -34 237581
rect 34 237547 46 237581
rect -46 237541 46 237547
rect -46 237473 46 237479
rect -46 237439 -34 237473
rect 34 237439 46 237473
rect -46 237433 46 237439
rect -102 237389 -56 237401
rect -102 236413 -96 237389
rect -62 236413 -56 237389
rect -102 236401 -56 236413
rect 56 237389 102 237401
rect 56 236413 62 237389
rect 96 236413 102 237389
rect 56 236401 102 236413
rect -46 236363 46 236369
rect -46 236329 -34 236363
rect 34 236329 46 236363
rect -46 236323 46 236329
rect -46 236255 46 236261
rect -46 236221 -34 236255
rect 34 236221 46 236255
rect -46 236215 46 236221
rect -102 236171 -56 236183
rect -102 235195 -96 236171
rect -62 235195 -56 236171
rect -102 235183 -56 235195
rect 56 236171 102 236183
rect 56 235195 62 236171
rect 96 235195 102 236171
rect 56 235183 102 235195
rect -46 235145 46 235151
rect -46 235111 -34 235145
rect 34 235111 46 235145
rect -46 235105 46 235111
rect -46 235037 46 235043
rect -46 235003 -34 235037
rect 34 235003 46 235037
rect -46 234997 46 235003
rect -102 234953 -56 234965
rect -102 233977 -96 234953
rect -62 233977 -56 234953
rect -102 233965 -56 233977
rect 56 234953 102 234965
rect 56 233977 62 234953
rect 96 233977 102 234953
rect 56 233965 102 233977
rect -46 233927 46 233933
rect -46 233893 -34 233927
rect 34 233893 46 233927
rect -46 233887 46 233893
rect -46 233819 46 233825
rect -46 233785 -34 233819
rect 34 233785 46 233819
rect -46 233779 46 233785
rect -102 233735 -56 233747
rect -102 232759 -96 233735
rect -62 232759 -56 233735
rect -102 232747 -56 232759
rect 56 233735 102 233747
rect 56 232759 62 233735
rect 96 232759 102 233735
rect 56 232747 102 232759
rect -46 232709 46 232715
rect -46 232675 -34 232709
rect 34 232675 46 232709
rect -46 232669 46 232675
rect -46 232601 46 232607
rect -46 232567 -34 232601
rect 34 232567 46 232601
rect -46 232561 46 232567
rect -102 232517 -56 232529
rect -102 231541 -96 232517
rect -62 231541 -56 232517
rect -102 231529 -56 231541
rect 56 232517 102 232529
rect 56 231541 62 232517
rect 96 231541 102 232517
rect 56 231529 102 231541
rect -46 231491 46 231497
rect -46 231457 -34 231491
rect 34 231457 46 231491
rect -46 231451 46 231457
rect -46 231383 46 231389
rect -46 231349 -34 231383
rect 34 231349 46 231383
rect -46 231343 46 231349
rect -102 231299 -56 231311
rect -102 230323 -96 231299
rect -62 230323 -56 231299
rect -102 230311 -56 230323
rect 56 231299 102 231311
rect 56 230323 62 231299
rect 96 230323 102 231299
rect 56 230311 102 230323
rect -46 230273 46 230279
rect -46 230239 -34 230273
rect 34 230239 46 230273
rect -46 230233 46 230239
rect -46 230165 46 230171
rect -46 230131 -34 230165
rect 34 230131 46 230165
rect -46 230125 46 230131
rect -102 230081 -56 230093
rect -102 229105 -96 230081
rect -62 229105 -56 230081
rect -102 229093 -56 229105
rect 56 230081 102 230093
rect 56 229105 62 230081
rect 96 229105 102 230081
rect 56 229093 102 229105
rect -46 229055 46 229061
rect -46 229021 -34 229055
rect 34 229021 46 229055
rect -46 229015 46 229021
rect -46 228947 46 228953
rect -46 228913 -34 228947
rect 34 228913 46 228947
rect -46 228907 46 228913
rect -102 228863 -56 228875
rect -102 227887 -96 228863
rect -62 227887 -56 228863
rect -102 227875 -56 227887
rect 56 228863 102 228875
rect 56 227887 62 228863
rect 96 227887 102 228863
rect 56 227875 102 227887
rect -46 227837 46 227843
rect -46 227803 -34 227837
rect 34 227803 46 227837
rect -46 227797 46 227803
rect -46 227729 46 227735
rect -46 227695 -34 227729
rect 34 227695 46 227729
rect -46 227689 46 227695
rect -102 227645 -56 227657
rect -102 226669 -96 227645
rect -62 226669 -56 227645
rect -102 226657 -56 226669
rect 56 227645 102 227657
rect 56 226669 62 227645
rect 96 226669 102 227645
rect 56 226657 102 226669
rect -46 226619 46 226625
rect -46 226585 -34 226619
rect 34 226585 46 226619
rect -46 226579 46 226585
rect -46 226511 46 226517
rect -46 226477 -34 226511
rect 34 226477 46 226511
rect -46 226471 46 226477
rect -102 226427 -56 226439
rect -102 225451 -96 226427
rect -62 225451 -56 226427
rect -102 225439 -56 225451
rect 56 226427 102 226439
rect 56 225451 62 226427
rect 96 225451 102 226427
rect 56 225439 102 225451
rect -46 225401 46 225407
rect -46 225367 -34 225401
rect 34 225367 46 225401
rect -46 225361 46 225367
rect -46 225293 46 225299
rect -46 225259 -34 225293
rect 34 225259 46 225293
rect -46 225253 46 225259
rect -102 225209 -56 225221
rect -102 224233 -96 225209
rect -62 224233 -56 225209
rect -102 224221 -56 224233
rect 56 225209 102 225221
rect 56 224233 62 225209
rect 96 224233 102 225209
rect 56 224221 102 224233
rect -46 224183 46 224189
rect -46 224149 -34 224183
rect 34 224149 46 224183
rect -46 224143 46 224149
rect -46 224075 46 224081
rect -46 224041 -34 224075
rect 34 224041 46 224075
rect -46 224035 46 224041
rect -102 223991 -56 224003
rect -102 223015 -96 223991
rect -62 223015 -56 223991
rect -102 223003 -56 223015
rect 56 223991 102 224003
rect 56 223015 62 223991
rect 96 223015 102 223991
rect 56 223003 102 223015
rect -46 222965 46 222971
rect -46 222931 -34 222965
rect 34 222931 46 222965
rect -46 222925 46 222931
rect -46 222857 46 222863
rect -46 222823 -34 222857
rect 34 222823 46 222857
rect -46 222817 46 222823
rect -102 222773 -56 222785
rect -102 221797 -96 222773
rect -62 221797 -56 222773
rect -102 221785 -56 221797
rect 56 222773 102 222785
rect 56 221797 62 222773
rect 96 221797 102 222773
rect 56 221785 102 221797
rect -46 221747 46 221753
rect -46 221713 -34 221747
rect 34 221713 46 221747
rect -46 221707 46 221713
rect -46 221639 46 221645
rect -46 221605 -34 221639
rect 34 221605 46 221639
rect -46 221599 46 221605
rect -102 221555 -56 221567
rect -102 220579 -96 221555
rect -62 220579 -56 221555
rect -102 220567 -56 220579
rect 56 221555 102 221567
rect 56 220579 62 221555
rect 96 220579 102 221555
rect 56 220567 102 220579
rect -46 220529 46 220535
rect -46 220495 -34 220529
rect 34 220495 46 220529
rect -46 220489 46 220495
rect -46 220421 46 220427
rect -46 220387 -34 220421
rect 34 220387 46 220421
rect -46 220381 46 220387
rect -102 220337 -56 220349
rect -102 219361 -96 220337
rect -62 219361 -56 220337
rect -102 219349 -56 219361
rect 56 220337 102 220349
rect 56 219361 62 220337
rect 96 219361 102 220337
rect 56 219349 102 219361
rect -46 219311 46 219317
rect -46 219277 -34 219311
rect 34 219277 46 219311
rect -46 219271 46 219277
rect -46 219203 46 219209
rect -46 219169 -34 219203
rect 34 219169 46 219203
rect -46 219163 46 219169
rect -102 219119 -56 219131
rect -102 218143 -96 219119
rect -62 218143 -56 219119
rect -102 218131 -56 218143
rect 56 219119 102 219131
rect 56 218143 62 219119
rect 96 218143 102 219119
rect 56 218131 102 218143
rect -46 218093 46 218099
rect -46 218059 -34 218093
rect 34 218059 46 218093
rect -46 218053 46 218059
rect -46 217985 46 217991
rect -46 217951 -34 217985
rect 34 217951 46 217985
rect -46 217945 46 217951
rect -102 217901 -56 217913
rect -102 216925 -96 217901
rect -62 216925 -56 217901
rect -102 216913 -56 216925
rect 56 217901 102 217913
rect 56 216925 62 217901
rect 96 216925 102 217901
rect 56 216913 102 216925
rect -46 216875 46 216881
rect -46 216841 -34 216875
rect 34 216841 46 216875
rect -46 216835 46 216841
rect -46 216767 46 216773
rect -46 216733 -34 216767
rect 34 216733 46 216767
rect -46 216727 46 216733
rect -102 216683 -56 216695
rect -102 215707 -96 216683
rect -62 215707 -56 216683
rect -102 215695 -56 215707
rect 56 216683 102 216695
rect 56 215707 62 216683
rect 96 215707 102 216683
rect 56 215695 102 215707
rect -46 215657 46 215663
rect -46 215623 -34 215657
rect 34 215623 46 215657
rect -46 215617 46 215623
rect -46 215549 46 215555
rect -46 215515 -34 215549
rect 34 215515 46 215549
rect -46 215509 46 215515
rect -102 215465 -56 215477
rect -102 214489 -96 215465
rect -62 214489 -56 215465
rect -102 214477 -56 214489
rect 56 215465 102 215477
rect 56 214489 62 215465
rect 96 214489 102 215465
rect 56 214477 102 214489
rect -46 214439 46 214445
rect -46 214405 -34 214439
rect 34 214405 46 214439
rect -46 214399 46 214405
rect -46 214331 46 214337
rect -46 214297 -34 214331
rect 34 214297 46 214331
rect -46 214291 46 214297
rect -102 214247 -56 214259
rect -102 213271 -96 214247
rect -62 213271 -56 214247
rect -102 213259 -56 213271
rect 56 214247 102 214259
rect 56 213271 62 214247
rect 96 213271 102 214247
rect 56 213259 102 213271
rect -46 213221 46 213227
rect -46 213187 -34 213221
rect 34 213187 46 213221
rect -46 213181 46 213187
rect -46 213113 46 213119
rect -46 213079 -34 213113
rect 34 213079 46 213113
rect -46 213073 46 213079
rect -102 213029 -56 213041
rect -102 212053 -96 213029
rect -62 212053 -56 213029
rect -102 212041 -56 212053
rect 56 213029 102 213041
rect 56 212053 62 213029
rect 96 212053 102 213029
rect 56 212041 102 212053
rect -46 212003 46 212009
rect -46 211969 -34 212003
rect 34 211969 46 212003
rect -46 211963 46 211969
rect -46 211895 46 211901
rect -46 211861 -34 211895
rect 34 211861 46 211895
rect -46 211855 46 211861
rect -102 211811 -56 211823
rect -102 210835 -96 211811
rect -62 210835 -56 211811
rect -102 210823 -56 210835
rect 56 211811 102 211823
rect 56 210835 62 211811
rect 96 210835 102 211811
rect 56 210823 102 210835
rect -46 210785 46 210791
rect -46 210751 -34 210785
rect 34 210751 46 210785
rect -46 210745 46 210751
rect -46 210677 46 210683
rect -46 210643 -34 210677
rect 34 210643 46 210677
rect -46 210637 46 210643
rect -102 210593 -56 210605
rect -102 209617 -96 210593
rect -62 209617 -56 210593
rect -102 209605 -56 209617
rect 56 210593 102 210605
rect 56 209617 62 210593
rect 96 209617 102 210593
rect 56 209605 102 209617
rect -46 209567 46 209573
rect -46 209533 -34 209567
rect 34 209533 46 209567
rect -46 209527 46 209533
rect -46 209459 46 209465
rect -46 209425 -34 209459
rect 34 209425 46 209459
rect -46 209419 46 209425
rect -102 209375 -56 209387
rect -102 208399 -96 209375
rect -62 208399 -56 209375
rect -102 208387 -56 208399
rect 56 209375 102 209387
rect 56 208399 62 209375
rect 96 208399 102 209375
rect 56 208387 102 208399
rect -46 208349 46 208355
rect -46 208315 -34 208349
rect 34 208315 46 208349
rect -46 208309 46 208315
rect -46 208241 46 208247
rect -46 208207 -34 208241
rect 34 208207 46 208241
rect -46 208201 46 208207
rect -102 208157 -56 208169
rect -102 207181 -96 208157
rect -62 207181 -56 208157
rect -102 207169 -56 207181
rect 56 208157 102 208169
rect 56 207181 62 208157
rect 96 207181 102 208157
rect 56 207169 102 207181
rect -46 207131 46 207137
rect -46 207097 -34 207131
rect 34 207097 46 207131
rect -46 207091 46 207097
rect -46 207023 46 207029
rect -46 206989 -34 207023
rect 34 206989 46 207023
rect -46 206983 46 206989
rect -102 206939 -56 206951
rect -102 205963 -96 206939
rect -62 205963 -56 206939
rect -102 205951 -56 205963
rect 56 206939 102 206951
rect 56 205963 62 206939
rect 96 205963 102 206939
rect 56 205951 102 205963
rect -46 205913 46 205919
rect -46 205879 -34 205913
rect 34 205879 46 205913
rect -46 205873 46 205879
rect -46 205805 46 205811
rect -46 205771 -34 205805
rect 34 205771 46 205805
rect -46 205765 46 205771
rect -102 205721 -56 205733
rect -102 204745 -96 205721
rect -62 204745 -56 205721
rect -102 204733 -56 204745
rect 56 205721 102 205733
rect 56 204745 62 205721
rect 96 204745 102 205721
rect 56 204733 102 204745
rect -46 204695 46 204701
rect -46 204661 -34 204695
rect 34 204661 46 204695
rect -46 204655 46 204661
rect -46 204587 46 204593
rect -46 204553 -34 204587
rect 34 204553 46 204587
rect -46 204547 46 204553
rect -102 204503 -56 204515
rect -102 203527 -96 204503
rect -62 203527 -56 204503
rect -102 203515 -56 203527
rect 56 204503 102 204515
rect 56 203527 62 204503
rect 96 203527 102 204503
rect 56 203515 102 203527
rect -46 203477 46 203483
rect -46 203443 -34 203477
rect 34 203443 46 203477
rect -46 203437 46 203443
rect -46 203369 46 203375
rect -46 203335 -34 203369
rect 34 203335 46 203369
rect -46 203329 46 203335
rect -102 203285 -56 203297
rect -102 202309 -96 203285
rect -62 202309 -56 203285
rect -102 202297 -56 202309
rect 56 203285 102 203297
rect 56 202309 62 203285
rect 96 202309 102 203285
rect 56 202297 102 202309
rect -46 202259 46 202265
rect -46 202225 -34 202259
rect 34 202225 46 202259
rect -46 202219 46 202225
rect -46 202151 46 202157
rect -46 202117 -34 202151
rect 34 202117 46 202151
rect -46 202111 46 202117
rect -102 202067 -56 202079
rect -102 201091 -96 202067
rect -62 201091 -56 202067
rect -102 201079 -56 201091
rect 56 202067 102 202079
rect 56 201091 62 202067
rect 96 201091 102 202067
rect 56 201079 102 201091
rect -46 201041 46 201047
rect -46 201007 -34 201041
rect 34 201007 46 201041
rect -46 201001 46 201007
rect -46 200933 46 200939
rect -46 200899 -34 200933
rect 34 200899 46 200933
rect -46 200893 46 200899
rect -102 200849 -56 200861
rect -102 199873 -96 200849
rect -62 199873 -56 200849
rect -102 199861 -56 199873
rect 56 200849 102 200861
rect 56 199873 62 200849
rect 96 199873 102 200849
rect 56 199861 102 199873
rect -46 199823 46 199829
rect -46 199789 -34 199823
rect 34 199789 46 199823
rect -46 199783 46 199789
rect -46 199715 46 199721
rect -46 199681 -34 199715
rect 34 199681 46 199715
rect -46 199675 46 199681
rect -102 199631 -56 199643
rect -102 198655 -96 199631
rect -62 198655 -56 199631
rect -102 198643 -56 198655
rect 56 199631 102 199643
rect 56 198655 62 199631
rect 96 198655 102 199631
rect 56 198643 102 198655
rect -46 198605 46 198611
rect -46 198571 -34 198605
rect 34 198571 46 198605
rect -46 198565 46 198571
rect -46 198497 46 198503
rect -46 198463 -34 198497
rect 34 198463 46 198497
rect -46 198457 46 198463
rect -102 198413 -56 198425
rect -102 197437 -96 198413
rect -62 197437 -56 198413
rect -102 197425 -56 197437
rect 56 198413 102 198425
rect 56 197437 62 198413
rect 96 197437 102 198413
rect 56 197425 102 197437
rect -46 197387 46 197393
rect -46 197353 -34 197387
rect 34 197353 46 197387
rect -46 197347 46 197353
rect -46 197279 46 197285
rect -46 197245 -34 197279
rect 34 197245 46 197279
rect -46 197239 46 197245
rect -102 197195 -56 197207
rect -102 196219 -96 197195
rect -62 196219 -56 197195
rect -102 196207 -56 196219
rect 56 197195 102 197207
rect 56 196219 62 197195
rect 96 196219 102 197195
rect 56 196207 102 196219
rect -46 196169 46 196175
rect -46 196135 -34 196169
rect 34 196135 46 196169
rect -46 196129 46 196135
rect -46 196061 46 196067
rect -46 196027 -34 196061
rect 34 196027 46 196061
rect -46 196021 46 196027
rect -102 195977 -56 195989
rect -102 195001 -96 195977
rect -62 195001 -56 195977
rect -102 194989 -56 195001
rect 56 195977 102 195989
rect 56 195001 62 195977
rect 96 195001 102 195977
rect 56 194989 102 195001
rect -46 194951 46 194957
rect -46 194917 -34 194951
rect 34 194917 46 194951
rect -46 194911 46 194917
rect -46 194843 46 194849
rect -46 194809 -34 194843
rect 34 194809 46 194843
rect -46 194803 46 194809
rect -102 194759 -56 194771
rect -102 193783 -96 194759
rect -62 193783 -56 194759
rect -102 193771 -56 193783
rect 56 194759 102 194771
rect 56 193783 62 194759
rect 96 193783 102 194759
rect 56 193771 102 193783
rect -46 193733 46 193739
rect -46 193699 -34 193733
rect 34 193699 46 193733
rect -46 193693 46 193699
rect -46 193625 46 193631
rect -46 193591 -34 193625
rect 34 193591 46 193625
rect -46 193585 46 193591
rect -102 193541 -56 193553
rect -102 192565 -96 193541
rect -62 192565 -56 193541
rect -102 192553 -56 192565
rect 56 193541 102 193553
rect 56 192565 62 193541
rect 96 192565 102 193541
rect 56 192553 102 192565
rect -46 192515 46 192521
rect -46 192481 -34 192515
rect 34 192481 46 192515
rect -46 192475 46 192481
rect -46 192407 46 192413
rect -46 192373 -34 192407
rect 34 192373 46 192407
rect -46 192367 46 192373
rect -102 192323 -56 192335
rect -102 191347 -96 192323
rect -62 191347 -56 192323
rect -102 191335 -56 191347
rect 56 192323 102 192335
rect 56 191347 62 192323
rect 96 191347 102 192323
rect 56 191335 102 191347
rect -46 191297 46 191303
rect -46 191263 -34 191297
rect 34 191263 46 191297
rect -46 191257 46 191263
rect -46 191189 46 191195
rect -46 191155 -34 191189
rect 34 191155 46 191189
rect -46 191149 46 191155
rect -102 191105 -56 191117
rect -102 190129 -96 191105
rect -62 190129 -56 191105
rect -102 190117 -56 190129
rect 56 191105 102 191117
rect 56 190129 62 191105
rect 96 190129 102 191105
rect 56 190117 102 190129
rect -46 190079 46 190085
rect -46 190045 -34 190079
rect 34 190045 46 190079
rect -46 190039 46 190045
rect -46 189971 46 189977
rect -46 189937 -34 189971
rect 34 189937 46 189971
rect -46 189931 46 189937
rect -102 189887 -56 189899
rect -102 188911 -96 189887
rect -62 188911 -56 189887
rect -102 188899 -56 188911
rect 56 189887 102 189899
rect 56 188911 62 189887
rect 96 188911 102 189887
rect 56 188899 102 188911
rect -46 188861 46 188867
rect -46 188827 -34 188861
rect 34 188827 46 188861
rect -46 188821 46 188827
rect -46 188753 46 188759
rect -46 188719 -34 188753
rect 34 188719 46 188753
rect -46 188713 46 188719
rect -102 188669 -56 188681
rect -102 187693 -96 188669
rect -62 187693 -56 188669
rect -102 187681 -56 187693
rect 56 188669 102 188681
rect 56 187693 62 188669
rect 96 187693 102 188669
rect 56 187681 102 187693
rect -46 187643 46 187649
rect -46 187609 -34 187643
rect 34 187609 46 187643
rect -46 187603 46 187609
rect -46 187535 46 187541
rect -46 187501 -34 187535
rect 34 187501 46 187535
rect -46 187495 46 187501
rect -102 187451 -56 187463
rect -102 186475 -96 187451
rect -62 186475 -56 187451
rect -102 186463 -56 186475
rect 56 187451 102 187463
rect 56 186475 62 187451
rect 96 186475 102 187451
rect 56 186463 102 186475
rect -46 186425 46 186431
rect -46 186391 -34 186425
rect 34 186391 46 186425
rect -46 186385 46 186391
rect -46 186317 46 186323
rect -46 186283 -34 186317
rect 34 186283 46 186317
rect -46 186277 46 186283
rect -102 186233 -56 186245
rect -102 185257 -96 186233
rect -62 185257 -56 186233
rect -102 185245 -56 185257
rect 56 186233 102 186245
rect 56 185257 62 186233
rect 96 185257 102 186233
rect 56 185245 102 185257
rect -46 185207 46 185213
rect -46 185173 -34 185207
rect 34 185173 46 185207
rect -46 185167 46 185173
rect -46 185099 46 185105
rect -46 185065 -34 185099
rect 34 185065 46 185099
rect -46 185059 46 185065
rect -102 185015 -56 185027
rect -102 184039 -96 185015
rect -62 184039 -56 185015
rect -102 184027 -56 184039
rect 56 185015 102 185027
rect 56 184039 62 185015
rect 96 184039 102 185015
rect 56 184027 102 184039
rect -46 183989 46 183995
rect -46 183955 -34 183989
rect 34 183955 46 183989
rect -46 183949 46 183955
rect -46 183881 46 183887
rect -46 183847 -34 183881
rect 34 183847 46 183881
rect -46 183841 46 183847
rect -102 183797 -56 183809
rect -102 182821 -96 183797
rect -62 182821 -56 183797
rect -102 182809 -56 182821
rect 56 183797 102 183809
rect 56 182821 62 183797
rect 96 182821 102 183797
rect 56 182809 102 182821
rect -46 182771 46 182777
rect -46 182737 -34 182771
rect 34 182737 46 182771
rect -46 182731 46 182737
rect -46 182663 46 182669
rect -46 182629 -34 182663
rect 34 182629 46 182663
rect -46 182623 46 182629
rect -102 182579 -56 182591
rect -102 181603 -96 182579
rect -62 181603 -56 182579
rect -102 181591 -56 181603
rect 56 182579 102 182591
rect 56 181603 62 182579
rect 96 181603 102 182579
rect 56 181591 102 181603
rect -46 181553 46 181559
rect -46 181519 -34 181553
rect 34 181519 46 181553
rect -46 181513 46 181519
rect -46 181445 46 181451
rect -46 181411 -34 181445
rect 34 181411 46 181445
rect -46 181405 46 181411
rect -102 181361 -56 181373
rect -102 180385 -96 181361
rect -62 180385 -56 181361
rect -102 180373 -56 180385
rect 56 181361 102 181373
rect 56 180385 62 181361
rect 96 180385 102 181361
rect 56 180373 102 180385
rect -46 180335 46 180341
rect -46 180301 -34 180335
rect 34 180301 46 180335
rect -46 180295 46 180301
rect -46 180227 46 180233
rect -46 180193 -34 180227
rect 34 180193 46 180227
rect -46 180187 46 180193
rect -102 180143 -56 180155
rect -102 179167 -96 180143
rect -62 179167 -56 180143
rect -102 179155 -56 179167
rect 56 180143 102 180155
rect 56 179167 62 180143
rect 96 179167 102 180143
rect 56 179155 102 179167
rect -46 179117 46 179123
rect -46 179083 -34 179117
rect 34 179083 46 179117
rect -46 179077 46 179083
rect -46 179009 46 179015
rect -46 178975 -34 179009
rect 34 178975 46 179009
rect -46 178969 46 178975
rect -102 178925 -56 178937
rect -102 177949 -96 178925
rect -62 177949 -56 178925
rect -102 177937 -56 177949
rect 56 178925 102 178937
rect 56 177949 62 178925
rect 96 177949 102 178925
rect 56 177937 102 177949
rect -46 177899 46 177905
rect -46 177865 -34 177899
rect 34 177865 46 177899
rect -46 177859 46 177865
rect -46 177791 46 177797
rect -46 177757 -34 177791
rect 34 177757 46 177791
rect -46 177751 46 177757
rect -102 177707 -56 177719
rect -102 176731 -96 177707
rect -62 176731 -56 177707
rect -102 176719 -56 176731
rect 56 177707 102 177719
rect 56 176731 62 177707
rect 96 176731 102 177707
rect 56 176719 102 176731
rect -46 176681 46 176687
rect -46 176647 -34 176681
rect 34 176647 46 176681
rect -46 176641 46 176647
rect -46 176573 46 176579
rect -46 176539 -34 176573
rect 34 176539 46 176573
rect -46 176533 46 176539
rect -102 176489 -56 176501
rect -102 175513 -96 176489
rect -62 175513 -56 176489
rect -102 175501 -56 175513
rect 56 176489 102 176501
rect 56 175513 62 176489
rect 96 175513 102 176489
rect 56 175501 102 175513
rect -46 175463 46 175469
rect -46 175429 -34 175463
rect 34 175429 46 175463
rect -46 175423 46 175429
rect -46 175355 46 175361
rect -46 175321 -34 175355
rect 34 175321 46 175355
rect -46 175315 46 175321
rect -102 175271 -56 175283
rect -102 174295 -96 175271
rect -62 174295 -56 175271
rect -102 174283 -56 174295
rect 56 175271 102 175283
rect 56 174295 62 175271
rect 96 174295 102 175271
rect 56 174283 102 174295
rect -46 174245 46 174251
rect -46 174211 -34 174245
rect 34 174211 46 174245
rect -46 174205 46 174211
rect -46 174137 46 174143
rect -46 174103 -34 174137
rect 34 174103 46 174137
rect -46 174097 46 174103
rect -102 174053 -56 174065
rect -102 173077 -96 174053
rect -62 173077 -56 174053
rect -102 173065 -56 173077
rect 56 174053 102 174065
rect 56 173077 62 174053
rect 96 173077 102 174053
rect 56 173065 102 173077
rect -46 173027 46 173033
rect -46 172993 -34 173027
rect 34 172993 46 173027
rect -46 172987 46 172993
rect -46 172919 46 172925
rect -46 172885 -34 172919
rect 34 172885 46 172919
rect -46 172879 46 172885
rect -102 172835 -56 172847
rect -102 171859 -96 172835
rect -62 171859 -56 172835
rect -102 171847 -56 171859
rect 56 172835 102 172847
rect 56 171859 62 172835
rect 96 171859 102 172835
rect 56 171847 102 171859
rect -46 171809 46 171815
rect -46 171775 -34 171809
rect 34 171775 46 171809
rect -46 171769 46 171775
rect -46 171701 46 171707
rect -46 171667 -34 171701
rect 34 171667 46 171701
rect -46 171661 46 171667
rect -102 171617 -56 171629
rect -102 170641 -96 171617
rect -62 170641 -56 171617
rect -102 170629 -56 170641
rect 56 171617 102 171629
rect 56 170641 62 171617
rect 96 170641 102 171617
rect 56 170629 102 170641
rect -46 170591 46 170597
rect -46 170557 -34 170591
rect 34 170557 46 170591
rect -46 170551 46 170557
rect -46 170483 46 170489
rect -46 170449 -34 170483
rect 34 170449 46 170483
rect -46 170443 46 170449
rect -102 170399 -56 170411
rect -102 169423 -96 170399
rect -62 169423 -56 170399
rect -102 169411 -56 169423
rect 56 170399 102 170411
rect 56 169423 62 170399
rect 96 169423 102 170399
rect 56 169411 102 169423
rect -46 169373 46 169379
rect -46 169339 -34 169373
rect 34 169339 46 169373
rect -46 169333 46 169339
rect -46 169265 46 169271
rect -46 169231 -34 169265
rect 34 169231 46 169265
rect -46 169225 46 169231
rect -102 169181 -56 169193
rect -102 168205 -96 169181
rect -62 168205 -56 169181
rect -102 168193 -56 168205
rect 56 169181 102 169193
rect 56 168205 62 169181
rect 96 168205 102 169181
rect 56 168193 102 168205
rect -46 168155 46 168161
rect -46 168121 -34 168155
rect 34 168121 46 168155
rect -46 168115 46 168121
rect -46 168047 46 168053
rect -46 168013 -34 168047
rect 34 168013 46 168047
rect -46 168007 46 168013
rect -102 167963 -56 167975
rect -102 166987 -96 167963
rect -62 166987 -56 167963
rect -102 166975 -56 166987
rect 56 167963 102 167975
rect 56 166987 62 167963
rect 96 166987 102 167963
rect 56 166975 102 166987
rect -46 166937 46 166943
rect -46 166903 -34 166937
rect 34 166903 46 166937
rect -46 166897 46 166903
rect -46 166829 46 166835
rect -46 166795 -34 166829
rect 34 166795 46 166829
rect -46 166789 46 166795
rect -102 166745 -56 166757
rect -102 165769 -96 166745
rect -62 165769 -56 166745
rect -102 165757 -56 165769
rect 56 166745 102 166757
rect 56 165769 62 166745
rect 96 165769 102 166745
rect 56 165757 102 165769
rect -46 165719 46 165725
rect -46 165685 -34 165719
rect 34 165685 46 165719
rect -46 165679 46 165685
rect -46 165611 46 165617
rect -46 165577 -34 165611
rect 34 165577 46 165611
rect -46 165571 46 165577
rect -102 165527 -56 165539
rect -102 164551 -96 165527
rect -62 164551 -56 165527
rect -102 164539 -56 164551
rect 56 165527 102 165539
rect 56 164551 62 165527
rect 96 164551 102 165527
rect 56 164539 102 164551
rect -46 164501 46 164507
rect -46 164467 -34 164501
rect 34 164467 46 164501
rect -46 164461 46 164467
rect -46 164393 46 164399
rect -46 164359 -34 164393
rect 34 164359 46 164393
rect -46 164353 46 164359
rect -102 164309 -56 164321
rect -102 163333 -96 164309
rect -62 163333 -56 164309
rect -102 163321 -56 163333
rect 56 164309 102 164321
rect 56 163333 62 164309
rect 96 163333 102 164309
rect 56 163321 102 163333
rect -46 163283 46 163289
rect -46 163249 -34 163283
rect 34 163249 46 163283
rect -46 163243 46 163249
rect -46 163175 46 163181
rect -46 163141 -34 163175
rect 34 163141 46 163175
rect -46 163135 46 163141
rect -102 163091 -56 163103
rect -102 162115 -96 163091
rect -62 162115 -56 163091
rect -102 162103 -56 162115
rect 56 163091 102 163103
rect 56 162115 62 163091
rect 96 162115 102 163091
rect 56 162103 102 162115
rect -46 162065 46 162071
rect -46 162031 -34 162065
rect 34 162031 46 162065
rect -46 162025 46 162031
rect -46 161957 46 161963
rect -46 161923 -34 161957
rect 34 161923 46 161957
rect -46 161917 46 161923
rect -102 161873 -56 161885
rect -102 160897 -96 161873
rect -62 160897 -56 161873
rect -102 160885 -56 160897
rect 56 161873 102 161885
rect 56 160897 62 161873
rect 96 160897 102 161873
rect 56 160885 102 160897
rect -46 160847 46 160853
rect -46 160813 -34 160847
rect 34 160813 46 160847
rect -46 160807 46 160813
rect -46 160739 46 160745
rect -46 160705 -34 160739
rect 34 160705 46 160739
rect -46 160699 46 160705
rect -102 160655 -56 160667
rect -102 159679 -96 160655
rect -62 159679 -56 160655
rect -102 159667 -56 159679
rect 56 160655 102 160667
rect 56 159679 62 160655
rect 96 159679 102 160655
rect 56 159667 102 159679
rect -46 159629 46 159635
rect -46 159595 -34 159629
rect 34 159595 46 159629
rect -46 159589 46 159595
rect -46 159521 46 159527
rect -46 159487 -34 159521
rect 34 159487 46 159521
rect -46 159481 46 159487
rect -102 159437 -56 159449
rect -102 158461 -96 159437
rect -62 158461 -56 159437
rect -102 158449 -56 158461
rect 56 159437 102 159449
rect 56 158461 62 159437
rect 96 158461 102 159437
rect 56 158449 102 158461
rect -46 158411 46 158417
rect -46 158377 -34 158411
rect 34 158377 46 158411
rect -46 158371 46 158377
rect -46 158303 46 158309
rect -46 158269 -34 158303
rect 34 158269 46 158303
rect -46 158263 46 158269
rect -102 158219 -56 158231
rect -102 157243 -96 158219
rect -62 157243 -56 158219
rect -102 157231 -56 157243
rect 56 158219 102 158231
rect 56 157243 62 158219
rect 96 157243 102 158219
rect 56 157231 102 157243
rect -46 157193 46 157199
rect -46 157159 -34 157193
rect 34 157159 46 157193
rect -46 157153 46 157159
rect -46 157085 46 157091
rect -46 157051 -34 157085
rect 34 157051 46 157085
rect -46 157045 46 157051
rect -102 157001 -56 157013
rect -102 156025 -96 157001
rect -62 156025 -56 157001
rect -102 156013 -56 156025
rect 56 157001 102 157013
rect 56 156025 62 157001
rect 96 156025 102 157001
rect 56 156013 102 156025
rect -46 155975 46 155981
rect -46 155941 -34 155975
rect 34 155941 46 155975
rect -46 155935 46 155941
rect -46 155867 46 155873
rect -46 155833 -34 155867
rect 34 155833 46 155867
rect -46 155827 46 155833
rect -102 155783 -56 155795
rect -102 154807 -96 155783
rect -62 154807 -56 155783
rect -102 154795 -56 154807
rect 56 155783 102 155795
rect 56 154807 62 155783
rect 96 154807 102 155783
rect 56 154795 102 154807
rect -46 154757 46 154763
rect -46 154723 -34 154757
rect 34 154723 46 154757
rect -46 154717 46 154723
rect -46 154649 46 154655
rect -46 154615 -34 154649
rect 34 154615 46 154649
rect -46 154609 46 154615
rect -102 154565 -56 154577
rect -102 153589 -96 154565
rect -62 153589 -56 154565
rect -102 153577 -56 153589
rect 56 154565 102 154577
rect 56 153589 62 154565
rect 96 153589 102 154565
rect 56 153577 102 153589
rect -46 153539 46 153545
rect -46 153505 -34 153539
rect 34 153505 46 153539
rect -46 153499 46 153505
rect -46 153431 46 153437
rect -46 153397 -34 153431
rect 34 153397 46 153431
rect -46 153391 46 153397
rect -102 153347 -56 153359
rect -102 152371 -96 153347
rect -62 152371 -56 153347
rect -102 152359 -56 152371
rect 56 153347 102 153359
rect 56 152371 62 153347
rect 96 152371 102 153347
rect 56 152359 102 152371
rect -46 152321 46 152327
rect -46 152287 -34 152321
rect 34 152287 46 152321
rect -46 152281 46 152287
rect -46 152213 46 152219
rect -46 152179 -34 152213
rect 34 152179 46 152213
rect -46 152173 46 152179
rect -102 152129 -56 152141
rect -102 151153 -96 152129
rect -62 151153 -56 152129
rect -102 151141 -56 151153
rect 56 152129 102 152141
rect 56 151153 62 152129
rect 96 151153 102 152129
rect 56 151141 102 151153
rect -46 151103 46 151109
rect -46 151069 -34 151103
rect 34 151069 46 151103
rect -46 151063 46 151069
rect -46 150995 46 151001
rect -46 150961 -34 150995
rect 34 150961 46 150995
rect -46 150955 46 150961
rect -102 150911 -56 150923
rect -102 149935 -96 150911
rect -62 149935 -56 150911
rect -102 149923 -56 149935
rect 56 150911 102 150923
rect 56 149935 62 150911
rect 96 149935 102 150911
rect 56 149923 102 149935
rect -46 149885 46 149891
rect -46 149851 -34 149885
rect 34 149851 46 149885
rect -46 149845 46 149851
rect -46 149777 46 149783
rect -46 149743 -34 149777
rect 34 149743 46 149777
rect -46 149737 46 149743
rect -102 149693 -56 149705
rect -102 148717 -96 149693
rect -62 148717 -56 149693
rect -102 148705 -56 148717
rect 56 149693 102 149705
rect 56 148717 62 149693
rect 96 148717 102 149693
rect 56 148705 102 148717
rect -46 148667 46 148673
rect -46 148633 -34 148667
rect 34 148633 46 148667
rect -46 148627 46 148633
rect -46 148559 46 148565
rect -46 148525 -34 148559
rect 34 148525 46 148559
rect -46 148519 46 148525
rect -102 148475 -56 148487
rect -102 147499 -96 148475
rect -62 147499 -56 148475
rect -102 147487 -56 147499
rect 56 148475 102 148487
rect 56 147499 62 148475
rect 96 147499 102 148475
rect 56 147487 102 147499
rect -46 147449 46 147455
rect -46 147415 -34 147449
rect 34 147415 46 147449
rect -46 147409 46 147415
rect -46 147341 46 147347
rect -46 147307 -34 147341
rect 34 147307 46 147341
rect -46 147301 46 147307
rect -102 147257 -56 147269
rect -102 146281 -96 147257
rect -62 146281 -56 147257
rect -102 146269 -56 146281
rect 56 147257 102 147269
rect 56 146281 62 147257
rect 96 146281 102 147257
rect 56 146269 102 146281
rect -46 146231 46 146237
rect -46 146197 -34 146231
rect 34 146197 46 146231
rect -46 146191 46 146197
rect -46 146123 46 146129
rect -46 146089 -34 146123
rect 34 146089 46 146123
rect -46 146083 46 146089
rect -102 146039 -56 146051
rect -102 145063 -96 146039
rect -62 145063 -56 146039
rect -102 145051 -56 145063
rect 56 146039 102 146051
rect 56 145063 62 146039
rect 96 145063 102 146039
rect 56 145051 102 145063
rect -46 145013 46 145019
rect -46 144979 -34 145013
rect 34 144979 46 145013
rect -46 144973 46 144979
rect -46 144905 46 144911
rect -46 144871 -34 144905
rect 34 144871 46 144905
rect -46 144865 46 144871
rect -102 144821 -56 144833
rect -102 143845 -96 144821
rect -62 143845 -56 144821
rect -102 143833 -56 143845
rect 56 144821 102 144833
rect 56 143845 62 144821
rect 96 143845 102 144821
rect 56 143833 102 143845
rect -46 143795 46 143801
rect -46 143761 -34 143795
rect 34 143761 46 143795
rect -46 143755 46 143761
rect -46 143687 46 143693
rect -46 143653 -34 143687
rect 34 143653 46 143687
rect -46 143647 46 143653
rect -102 143603 -56 143615
rect -102 142627 -96 143603
rect -62 142627 -56 143603
rect -102 142615 -56 142627
rect 56 143603 102 143615
rect 56 142627 62 143603
rect 96 142627 102 143603
rect 56 142615 102 142627
rect -46 142577 46 142583
rect -46 142543 -34 142577
rect 34 142543 46 142577
rect -46 142537 46 142543
rect -46 142469 46 142475
rect -46 142435 -34 142469
rect 34 142435 46 142469
rect -46 142429 46 142435
rect -102 142385 -56 142397
rect -102 141409 -96 142385
rect -62 141409 -56 142385
rect -102 141397 -56 141409
rect 56 142385 102 142397
rect 56 141409 62 142385
rect 96 141409 102 142385
rect 56 141397 102 141409
rect -46 141359 46 141365
rect -46 141325 -34 141359
rect 34 141325 46 141359
rect -46 141319 46 141325
rect -46 141251 46 141257
rect -46 141217 -34 141251
rect 34 141217 46 141251
rect -46 141211 46 141217
rect -102 141167 -56 141179
rect -102 140191 -96 141167
rect -62 140191 -56 141167
rect -102 140179 -56 140191
rect 56 141167 102 141179
rect 56 140191 62 141167
rect 96 140191 102 141167
rect 56 140179 102 140191
rect -46 140141 46 140147
rect -46 140107 -34 140141
rect 34 140107 46 140141
rect -46 140101 46 140107
rect -46 140033 46 140039
rect -46 139999 -34 140033
rect 34 139999 46 140033
rect -46 139993 46 139999
rect -102 139949 -56 139961
rect -102 138973 -96 139949
rect -62 138973 -56 139949
rect -102 138961 -56 138973
rect 56 139949 102 139961
rect 56 138973 62 139949
rect 96 138973 102 139949
rect 56 138961 102 138973
rect -46 138923 46 138929
rect -46 138889 -34 138923
rect 34 138889 46 138923
rect -46 138883 46 138889
rect -46 138815 46 138821
rect -46 138781 -34 138815
rect 34 138781 46 138815
rect -46 138775 46 138781
rect -102 138731 -56 138743
rect -102 137755 -96 138731
rect -62 137755 -56 138731
rect -102 137743 -56 137755
rect 56 138731 102 138743
rect 56 137755 62 138731
rect 96 137755 102 138731
rect 56 137743 102 137755
rect -46 137705 46 137711
rect -46 137671 -34 137705
rect 34 137671 46 137705
rect -46 137665 46 137671
rect -46 137597 46 137603
rect -46 137563 -34 137597
rect 34 137563 46 137597
rect -46 137557 46 137563
rect -102 137513 -56 137525
rect -102 136537 -96 137513
rect -62 136537 -56 137513
rect -102 136525 -56 136537
rect 56 137513 102 137525
rect 56 136537 62 137513
rect 96 136537 102 137513
rect 56 136525 102 136537
rect -46 136487 46 136493
rect -46 136453 -34 136487
rect 34 136453 46 136487
rect -46 136447 46 136453
rect -46 136379 46 136385
rect -46 136345 -34 136379
rect 34 136345 46 136379
rect -46 136339 46 136345
rect -102 136295 -56 136307
rect -102 135319 -96 136295
rect -62 135319 -56 136295
rect -102 135307 -56 135319
rect 56 136295 102 136307
rect 56 135319 62 136295
rect 96 135319 102 136295
rect 56 135307 102 135319
rect -46 135269 46 135275
rect -46 135235 -34 135269
rect 34 135235 46 135269
rect -46 135229 46 135235
rect -46 135161 46 135167
rect -46 135127 -34 135161
rect 34 135127 46 135161
rect -46 135121 46 135127
rect -102 135077 -56 135089
rect -102 134101 -96 135077
rect -62 134101 -56 135077
rect -102 134089 -56 134101
rect 56 135077 102 135089
rect 56 134101 62 135077
rect 96 134101 102 135077
rect 56 134089 102 134101
rect -46 134051 46 134057
rect -46 134017 -34 134051
rect 34 134017 46 134051
rect -46 134011 46 134017
rect -46 133943 46 133949
rect -46 133909 -34 133943
rect 34 133909 46 133943
rect -46 133903 46 133909
rect -102 133859 -56 133871
rect -102 132883 -96 133859
rect -62 132883 -56 133859
rect -102 132871 -56 132883
rect 56 133859 102 133871
rect 56 132883 62 133859
rect 96 132883 102 133859
rect 56 132871 102 132883
rect -46 132833 46 132839
rect -46 132799 -34 132833
rect 34 132799 46 132833
rect -46 132793 46 132799
rect -46 132725 46 132731
rect -46 132691 -34 132725
rect 34 132691 46 132725
rect -46 132685 46 132691
rect -102 132641 -56 132653
rect -102 131665 -96 132641
rect -62 131665 -56 132641
rect -102 131653 -56 131665
rect 56 132641 102 132653
rect 56 131665 62 132641
rect 96 131665 102 132641
rect 56 131653 102 131665
rect -46 131615 46 131621
rect -46 131581 -34 131615
rect 34 131581 46 131615
rect -46 131575 46 131581
rect -46 131507 46 131513
rect -46 131473 -34 131507
rect 34 131473 46 131507
rect -46 131467 46 131473
rect -102 131423 -56 131435
rect -102 130447 -96 131423
rect -62 130447 -56 131423
rect -102 130435 -56 130447
rect 56 131423 102 131435
rect 56 130447 62 131423
rect 96 130447 102 131423
rect 56 130435 102 130447
rect -46 130397 46 130403
rect -46 130363 -34 130397
rect 34 130363 46 130397
rect -46 130357 46 130363
rect -46 130289 46 130295
rect -46 130255 -34 130289
rect 34 130255 46 130289
rect -46 130249 46 130255
rect -102 130205 -56 130217
rect -102 129229 -96 130205
rect -62 129229 -56 130205
rect -102 129217 -56 129229
rect 56 130205 102 130217
rect 56 129229 62 130205
rect 96 129229 102 130205
rect 56 129217 102 129229
rect -46 129179 46 129185
rect -46 129145 -34 129179
rect 34 129145 46 129179
rect -46 129139 46 129145
rect -46 129071 46 129077
rect -46 129037 -34 129071
rect 34 129037 46 129071
rect -46 129031 46 129037
rect -102 128987 -56 128999
rect -102 128011 -96 128987
rect -62 128011 -56 128987
rect -102 127999 -56 128011
rect 56 128987 102 128999
rect 56 128011 62 128987
rect 96 128011 102 128987
rect 56 127999 102 128011
rect -46 127961 46 127967
rect -46 127927 -34 127961
rect 34 127927 46 127961
rect -46 127921 46 127927
rect -46 127853 46 127859
rect -46 127819 -34 127853
rect 34 127819 46 127853
rect -46 127813 46 127819
rect -102 127769 -56 127781
rect -102 126793 -96 127769
rect -62 126793 -56 127769
rect -102 126781 -56 126793
rect 56 127769 102 127781
rect 56 126793 62 127769
rect 96 126793 102 127769
rect 56 126781 102 126793
rect -46 126743 46 126749
rect -46 126709 -34 126743
rect 34 126709 46 126743
rect -46 126703 46 126709
rect -46 126635 46 126641
rect -46 126601 -34 126635
rect 34 126601 46 126635
rect -46 126595 46 126601
rect -102 126551 -56 126563
rect -102 125575 -96 126551
rect -62 125575 -56 126551
rect -102 125563 -56 125575
rect 56 126551 102 126563
rect 56 125575 62 126551
rect 96 125575 102 126551
rect 56 125563 102 125575
rect -46 125525 46 125531
rect -46 125491 -34 125525
rect 34 125491 46 125525
rect -46 125485 46 125491
rect -46 125417 46 125423
rect -46 125383 -34 125417
rect 34 125383 46 125417
rect -46 125377 46 125383
rect -102 125333 -56 125345
rect -102 124357 -96 125333
rect -62 124357 -56 125333
rect -102 124345 -56 124357
rect 56 125333 102 125345
rect 56 124357 62 125333
rect 96 124357 102 125333
rect 56 124345 102 124357
rect -46 124307 46 124313
rect -46 124273 -34 124307
rect 34 124273 46 124307
rect -46 124267 46 124273
rect -46 124199 46 124205
rect -46 124165 -34 124199
rect 34 124165 46 124199
rect -46 124159 46 124165
rect -102 124115 -56 124127
rect -102 123139 -96 124115
rect -62 123139 -56 124115
rect -102 123127 -56 123139
rect 56 124115 102 124127
rect 56 123139 62 124115
rect 96 123139 102 124115
rect 56 123127 102 123139
rect -46 123089 46 123095
rect -46 123055 -34 123089
rect 34 123055 46 123089
rect -46 123049 46 123055
rect -46 122981 46 122987
rect -46 122947 -34 122981
rect 34 122947 46 122981
rect -46 122941 46 122947
rect -102 122897 -56 122909
rect -102 121921 -96 122897
rect -62 121921 -56 122897
rect -102 121909 -56 121921
rect 56 122897 102 122909
rect 56 121921 62 122897
rect 96 121921 102 122897
rect 56 121909 102 121921
rect -46 121871 46 121877
rect -46 121837 -34 121871
rect 34 121837 46 121871
rect -46 121831 46 121837
rect -46 121763 46 121769
rect -46 121729 -34 121763
rect 34 121729 46 121763
rect -46 121723 46 121729
rect -102 121679 -56 121691
rect -102 120703 -96 121679
rect -62 120703 -56 121679
rect -102 120691 -56 120703
rect 56 121679 102 121691
rect 56 120703 62 121679
rect 96 120703 102 121679
rect 56 120691 102 120703
rect -46 120653 46 120659
rect -46 120619 -34 120653
rect 34 120619 46 120653
rect -46 120613 46 120619
rect -46 120545 46 120551
rect -46 120511 -34 120545
rect 34 120511 46 120545
rect -46 120505 46 120511
rect -102 120461 -56 120473
rect -102 119485 -96 120461
rect -62 119485 -56 120461
rect -102 119473 -56 119485
rect 56 120461 102 120473
rect 56 119485 62 120461
rect 96 119485 102 120461
rect 56 119473 102 119485
rect -46 119435 46 119441
rect -46 119401 -34 119435
rect 34 119401 46 119435
rect -46 119395 46 119401
rect -46 119327 46 119333
rect -46 119293 -34 119327
rect 34 119293 46 119327
rect -46 119287 46 119293
rect -102 119243 -56 119255
rect -102 118267 -96 119243
rect -62 118267 -56 119243
rect -102 118255 -56 118267
rect 56 119243 102 119255
rect 56 118267 62 119243
rect 96 118267 102 119243
rect 56 118255 102 118267
rect -46 118217 46 118223
rect -46 118183 -34 118217
rect 34 118183 46 118217
rect -46 118177 46 118183
rect -46 118109 46 118115
rect -46 118075 -34 118109
rect 34 118075 46 118109
rect -46 118069 46 118075
rect -102 118025 -56 118037
rect -102 117049 -96 118025
rect -62 117049 -56 118025
rect -102 117037 -56 117049
rect 56 118025 102 118037
rect 56 117049 62 118025
rect 96 117049 102 118025
rect 56 117037 102 117049
rect -46 116999 46 117005
rect -46 116965 -34 116999
rect 34 116965 46 116999
rect -46 116959 46 116965
rect -46 116891 46 116897
rect -46 116857 -34 116891
rect 34 116857 46 116891
rect -46 116851 46 116857
rect -102 116807 -56 116819
rect -102 115831 -96 116807
rect -62 115831 -56 116807
rect -102 115819 -56 115831
rect 56 116807 102 116819
rect 56 115831 62 116807
rect 96 115831 102 116807
rect 56 115819 102 115831
rect -46 115781 46 115787
rect -46 115747 -34 115781
rect 34 115747 46 115781
rect -46 115741 46 115747
rect -46 115673 46 115679
rect -46 115639 -34 115673
rect 34 115639 46 115673
rect -46 115633 46 115639
rect -102 115589 -56 115601
rect -102 114613 -96 115589
rect -62 114613 -56 115589
rect -102 114601 -56 114613
rect 56 115589 102 115601
rect 56 114613 62 115589
rect 96 114613 102 115589
rect 56 114601 102 114613
rect -46 114563 46 114569
rect -46 114529 -34 114563
rect 34 114529 46 114563
rect -46 114523 46 114529
rect -46 114455 46 114461
rect -46 114421 -34 114455
rect 34 114421 46 114455
rect -46 114415 46 114421
rect -102 114371 -56 114383
rect -102 113395 -96 114371
rect -62 113395 -56 114371
rect -102 113383 -56 113395
rect 56 114371 102 114383
rect 56 113395 62 114371
rect 96 113395 102 114371
rect 56 113383 102 113395
rect -46 113345 46 113351
rect -46 113311 -34 113345
rect 34 113311 46 113345
rect -46 113305 46 113311
rect -46 113237 46 113243
rect -46 113203 -34 113237
rect 34 113203 46 113237
rect -46 113197 46 113203
rect -102 113153 -56 113165
rect -102 112177 -96 113153
rect -62 112177 -56 113153
rect -102 112165 -56 112177
rect 56 113153 102 113165
rect 56 112177 62 113153
rect 96 112177 102 113153
rect 56 112165 102 112177
rect -46 112127 46 112133
rect -46 112093 -34 112127
rect 34 112093 46 112127
rect -46 112087 46 112093
rect -46 112019 46 112025
rect -46 111985 -34 112019
rect 34 111985 46 112019
rect -46 111979 46 111985
rect -102 111935 -56 111947
rect -102 110959 -96 111935
rect -62 110959 -56 111935
rect -102 110947 -56 110959
rect 56 111935 102 111947
rect 56 110959 62 111935
rect 96 110959 102 111935
rect 56 110947 102 110959
rect -46 110909 46 110915
rect -46 110875 -34 110909
rect 34 110875 46 110909
rect -46 110869 46 110875
rect -46 110801 46 110807
rect -46 110767 -34 110801
rect 34 110767 46 110801
rect -46 110761 46 110767
rect -102 110717 -56 110729
rect -102 109741 -96 110717
rect -62 109741 -56 110717
rect -102 109729 -56 109741
rect 56 110717 102 110729
rect 56 109741 62 110717
rect 96 109741 102 110717
rect 56 109729 102 109741
rect -46 109691 46 109697
rect -46 109657 -34 109691
rect 34 109657 46 109691
rect -46 109651 46 109657
rect -46 109583 46 109589
rect -46 109549 -34 109583
rect 34 109549 46 109583
rect -46 109543 46 109549
rect -102 109499 -56 109511
rect -102 108523 -96 109499
rect -62 108523 -56 109499
rect -102 108511 -56 108523
rect 56 109499 102 109511
rect 56 108523 62 109499
rect 96 108523 102 109499
rect 56 108511 102 108523
rect -46 108473 46 108479
rect -46 108439 -34 108473
rect 34 108439 46 108473
rect -46 108433 46 108439
rect -46 108365 46 108371
rect -46 108331 -34 108365
rect 34 108331 46 108365
rect -46 108325 46 108331
rect -102 108281 -56 108293
rect -102 107305 -96 108281
rect -62 107305 -56 108281
rect -102 107293 -56 107305
rect 56 108281 102 108293
rect 56 107305 62 108281
rect 96 107305 102 108281
rect 56 107293 102 107305
rect -46 107255 46 107261
rect -46 107221 -34 107255
rect 34 107221 46 107255
rect -46 107215 46 107221
rect -46 107147 46 107153
rect -46 107113 -34 107147
rect 34 107113 46 107147
rect -46 107107 46 107113
rect -102 107063 -56 107075
rect -102 106087 -96 107063
rect -62 106087 -56 107063
rect -102 106075 -56 106087
rect 56 107063 102 107075
rect 56 106087 62 107063
rect 96 106087 102 107063
rect 56 106075 102 106087
rect -46 106037 46 106043
rect -46 106003 -34 106037
rect 34 106003 46 106037
rect -46 105997 46 106003
rect -46 105929 46 105935
rect -46 105895 -34 105929
rect 34 105895 46 105929
rect -46 105889 46 105895
rect -102 105845 -56 105857
rect -102 104869 -96 105845
rect -62 104869 -56 105845
rect -102 104857 -56 104869
rect 56 105845 102 105857
rect 56 104869 62 105845
rect 96 104869 102 105845
rect 56 104857 102 104869
rect -46 104819 46 104825
rect -46 104785 -34 104819
rect 34 104785 46 104819
rect -46 104779 46 104785
rect -46 104711 46 104717
rect -46 104677 -34 104711
rect 34 104677 46 104711
rect -46 104671 46 104677
rect -102 104627 -56 104639
rect -102 103651 -96 104627
rect -62 103651 -56 104627
rect -102 103639 -56 103651
rect 56 104627 102 104639
rect 56 103651 62 104627
rect 96 103651 102 104627
rect 56 103639 102 103651
rect -46 103601 46 103607
rect -46 103567 -34 103601
rect 34 103567 46 103601
rect -46 103561 46 103567
rect -46 103493 46 103499
rect -46 103459 -34 103493
rect 34 103459 46 103493
rect -46 103453 46 103459
rect -102 103409 -56 103421
rect -102 102433 -96 103409
rect -62 102433 -56 103409
rect -102 102421 -56 102433
rect 56 103409 102 103421
rect 56 102433 62 103409
rect 96 102433 102 103409
rect 56 102421 102 102433
rect -46 102383 46 102389
rect -46 102349 -34 102383
rect 34 102349 46 102383
rect -46 102343 46 102349
rect -46 102275 46 102281
rect -46 102241 -34 102275
rect 34 102241 46 102275
rect -46 102235 46 102241
rect -102 102191 -56 102203
rect -102 101215 -96 102191
rect -62 101215 -56 102191
rect -102 101203 -56 101215
rect 56 102191 102 102203
rect 56 101215 62 102191
rect 96 101215 102 102191
rect 56 101203 102 101215
rect -46 101165 46 101171
rect -46 101131 -34 101165
rect 34 101131 46 101165
rect -46 101125 46 101131
rect -46 101057 46 101063
rect -46 101023 -34 101057
rect 34 101023 46 101057
rect -46 101017 46 101023
rect -102 100973 -56 100985
rect -102 99997 -96 100973
rect -62 99997 -56 100973
rect -102 99985 -56 99997
rect 56 100973 102 100985
rect 56 99997 62 100973
rect 96 99997 102 100973
rect 56 99985 102 99997
rect -46 99947 46 99953
rect -46 99913 -34 99947
rect 34 99913 46 99947
rect -46 99907 46 99913
rect -46 99839 46 99845
rect -46 99805 -34 99839
rect 34 99805 46 99839
rect -46 99799 46 99805
rect -102 99755 -56 99767
rect -102 98779 -96 99755
rect -62 98779 -56 99755
rect -102 98767 -56 98779
rect 56 99755 102 99767
rect 56 98779 62 99755
rect 96 98779 102 99755
rect 56 98767 102 98779
rect -46 98729 46 98735
rect -46 98695 -34 98729
rect 34 98695 46 98729
rect -46 98689 46 98695
rect -46 98621 46 98627
rect -46 98587 -34 98621
rect 34 98587 46 98621
rect -46 98581 46 98587
rect -102 98537 -56 98549
rect -102 97561 -96 98537
rect -62 97561 -56 98537
rect -102 97549 -56 97561
rect 56 98537 102 98549
rect 56 97561 62 98537
rect 96 97561 102 98537
rect 56 97549 102 97561
rect -46 97511 46 97517
rect -46 97477 -34 97511
rect 34 97477 46 97511
rect -46 97471 46 97477
rect -46 97403 46 97409
rect -46 97369 -34 97403
rect 34 97369 46 97403
rect -46 97363 46 97369
rect -102 97319 -56 97331
rect -102 96343 -96 97319
rect -62 96343 -56 97319
rect -102 96331 -56 96343
rect 56 97319 102 97331
rect 56 96343 62 97319
rect 96 96343 102 97319
rect 56 96331 102 96343
rect -46 96293 46 96299
rect -46 96259 -34 96293
rect 34 96259 46 96293
rect -46 96253 46 96259
rect -46 96185 46 96191
rect -46 96151 -34 96185
rect 34 96151 46 96185
rect -46 96145 46 96151
rect -102 96101 -56 96113
rect -102 95125 -96 96101
rect -62 95125 -56 96101
rect -102 95113 -56 95125
rect 56 96101 102 96113
rect 56 95125 62 96101
rect 96 95125 102 96101
rect 56 95113 102 95125
rect -46 95075 46 95081
rect -46 95041 -34 95075
rect 34 95041 46 95075
rect -46 95035 46 95041
rect -46 94967 46 94973
rect -46 94933 -34 94967
rect 34 94933 46 94967
rect -46 94927 46 94933
rect -102 94883 -56 94895
rect -102 93907 -96 94883
rect -62 93907 -56 94883
rect -102 93895 -56 93907
rect 56 94883 102 94895
rect 56 93907 62 94883
rect 96 93907 102 94883
rect 56 93895 102 93907
rect -46 93857 46 93863
rect -46 93823 -34 93857
rect 34 93823 46 93857
rect -46 93817 46 93823
rect -46 93749 46 93755
rect -46 93715 -34 93749
rect 34 93715 46 93749
rect -46 93709 46 93715
rect -102 93665 -56 93677
rect -102 92689 -96 93665
rect -62 92689 -56 93665
rect -102 92677 -56 92689
rect 56 93665 102 93677
rect 56 92689 62 93665
rect 96 92689 102 93665
rect 56 92677 102 92689
rect -46 92639 46 92645
rect -46 92605 -34 92639
rect 34 92605 46 92639
rect -46 92599 46 92605
rect -46 92531 46 92537
rect -46 92497 -34 92531
rect 34 92497 46 92531
rect -46 92491 46 92497
rect -102 92447 -56 92459
rect -102 91471 -96 92447
rect -62 91471 -56 92447
rect -102 91459 -56 91471
rect 56 92447 102 92459
rect 56 91471 62 92447
rect 96 91471 102 92447
rect 56 91459 102 91471
rect -46 91421 46 91427
rect -46 91387 -34 91421
rect 34 91387 46 91421
rect -46 91381 46 91387
rect -46 91313 46 91319
rect -46 91279 -34 91313
rect 34 91279 46 91313
rect -46 91273 46 91279
rect -102 91229 -56 91241
rect -102 90253 -96 91229
rect -62 90253 -56 91229
rect -102 90241 -56 90253
rect 56 91229 102 91241
rect 56 90253 62 91229
rect 96 90253 102 91229
rect 56 90241 102 90253
rect -46 90203 46 90209
rect -46 90169 -34 90203
rect 34 90169 46 90203
rect -46 90163 46 90169
rect -46 90095 46 90101
rect -46 90061 -34 90095
rect 34 90061 46 90095
rect -46 90055 46 90061
rect -102 90011 -56 90023
rect -102 89035 -96 90011
rect -62 89035 -56 90011
rect -102 89023 -56 89035
rect 56 90011 102 90023
rect 56 89035 62 90011
rect 96 89035 102 90011
rect 56 89023 102 89035
rect -46 88985 46 88991
rect -46 88951 -34 88985
rect 34 88951 46 88985
rect -46 88945 46 88951
rect -46 88877 46 88883
rect -46 88843 -34 88877
rect 34 88843 46 88877
rect -46 88837 46 88843
rect -102 88793 -56 88805
rect -102 87817 -96 88793
rect -62 87817 -56 88793
rect -102 87805 -56 87817
rect 56 88793 102 88805
rect 56 87817 62 88793
rect 96 87817 102 88793
rect 56 87805 102 87817
rect -46 87767 46 87773
rect -46 87733 -34 87767
rect 34 87733 46 87767
rect -46 87727 46 87733
rect -46 87659 46 87665
rect -46 87625 -34 87659
rect 34 87625 46 87659
rect -46 87619 46 87625
rect -102 87575 -56 87587
rect -102 86599 -96 87575
rect -62 86599 -56 87575
rect -102 86587 -56 86599
rect 56 87575 102 87587
rect 56 86599 62 87575
rect 96 86599 102 87575
rect 56 86587 102 86599
rect -46 86549 46 86555
rect -46 86515 -34 86549
rect 34 86515 46 86549
rect -46 86509 46 86515
rect -46 86441 46 86447
rect -46 86407 -34 86441
rect 34 86407 46 86441
rect -46 86401 46 86407
rect -102 86357 -56 86369
rect -102 85381 -96 86357
rect -62 85381 -56 86357
rect -102 85369 -56 85381
rect 56 86357 102 86369
rect 56 85381 62 86357
rect 96 85381 102 86357
rect 56 85369 102 85381
rect -46 85331 46 85337
rect -46 85297 -34 85331
rect 34 85297 46 85331
rect -46 85291 46 85297
rect -46 85223 46 85229
rect -46 85189 -34 85223
rect 34 85189 46 85223
rect -46 85183 46 85189
rect -102 85139 -56 85151
rect -102 84163 -96 85139
rect -62 84163 -56 85139
rect -102 84151 -56 84163
rect 56 85139 102 85151
rect 56 84163 62 85139
rect 96 84163 102 85139
rect 56 84151 102 84163
rect -46 84113 46 84119
rect -46 84079 -34 84113
rect 34 84079 46 84113
rect -46 84073 46 84079
rect -46 84005 46 84011
rect -46 83971 -34 84005
rect 34 83971 46 84005
rect -46 83965 46 83971
rect -102 83921 -56 83933
rect -102 82945 -96 83921
rect -62 82945 -56 83921
rect -102 82933 -56 82945
rect 56 83921 102 83933
rect 56 82945 62 83921
rect 96 82945 102 83921
rect 56 82933 102 82945
rect -46 82895 46 82901
rect -46 82861 -34 82895
rect 34 82861 46 82895
rect -46 82855 46 82861
rect -46 82787 46 82793
rect -46 82753 -34 82787
rect 34 82753 46 82787
rect -46 82747 46 82753
rect -102 82703 -56 82715
rect -102 81727 -96 82703
rect -62 81727 -56 82703
rect -102 81715 -56 81727
rect 56 82703 102 82715
rect 56 81727 62 82703
rect 96 81727 102 82703
rect 56 81715 102 81727
rect -46 81677 46 81683
rect -46 81643 -34 81677
rect 34 81643 46 81677
rect -46 81637 46 81643
rect -46 81569 46 81575
rect -46 81535 -34 81569
rect 34 81535 46 81569
rect -46 81529 46 81535
rect -102 81485 -56 81497
rect -102 80509 -96 81485
rect -62 80509 -56 81485
rect -102 80497 -56 80509
rect 56 81485 102 81497
rect 56 80509 62 81485
rect 96 80509 102 81485
rect 56 80497 102 80509
rect -46 80459 46 80465
rect -46 80425 -34 80459
rect 34 80425 46 80459
rect -46 80419 46 80425
rect -46 80351 46 80357
rect -46 80317 -34 80351
rect 34 80317 46 80351
rect -46 80311 46 80317
rect -102 80267 -56 80279
rect -102 79291 -96 80267
rect -62 79291 -56 80267
rect -102 79279 -56 79291
rect 56 80267 102 80279
rect 56 79291 62 80267
rect 96 79291 102 80267
rect 56 79279 102 79291
rect -46 79241 46 79247
rect -46 79207 -34 79241
rect 34 79207 46 79241
rect -46 79201 46 79207
rect -46 79133 46 79139
rect -46 79099 -34 79133
rect 34 79099 46 79133
rect -46 79093 46 79099
rect -102 79049 -56 79061
rect -102 78073 -96 79049
rect -62 78073 -56 79049
rect -102 78061 -56 78073
rect 56 79049 102 79061
rect 56 78073 62 79049
rect 96 78073 102 79049
rect 56 78061 102 78073
rect -46 78023 46 78029
rect -46 77989 -34 78023
rect 34 77989 46 78023
rect -46 77983 46 77989
rect -46 77915 46 77921
rect -46 77881 -34 77915
rect 34 77881 46 77915
rect -46 77875 46 77881
rect -102 77831 -56 77843
rect -102 76855 -96 77831
rect -62 76855 -56 77831
rect -102 76843 -56 76855
rect 56 77831 102 77843
rect 56 76855 62 77831
rect 96 76855 102 77831
rect 56 76843 102 76855
rect -46 76805 46 76811
rect -46 76771 -34 76805
rect 34 76771 46 76805
rect -46 76765 46 76771
rect -46 76697 46 76703
rect -46 76663 -34 76697
rect 34 76663 46 76697
rect -46 76657 46 76663
rect -102 76613 -56 76625
rect -102 75637 -96 76613
rect -62 75637 -56 76613
rect -102 75625 -56 75637
rect 56 76613 102 76625
rect 56 75637 62 76613
rect 96 75637 102 76613
rect 56 75625 102 75637
rect -46 75587 46 75593
rect -46 75553 -34 75587
rect 34 75553 46 75587
rect -46 75547 46 75553
rect -46 75479 46 75485
rect -46 75445 -34 75479
rect 34 75445 46 75479
rect -46 75439 46 75445
rect -102 75395 -56 75407
rect -102 74419 -96 75395
rect -62 74419 -56 75395
rect -102 74407 -56 74419
rect 56 75395 102 75407
rect 56 74419 62 75395
rect 96 74419 102 75395
rect 56 74407 102 74419
rect -46 74369 46 74375
rect -46 74335 -34 74369
rect 34 74335 46 74369
rect -46 74329 46 74335
rect -46 74261 46 74267
rect -46 74227 -34 74261
rect 34 74227 46 74261
rect -46 74221 46 74227
rect -102 74177 -56 74189
rect -102 73201 -96 74177
rect -62 73201 -56 74177
rect -102 73189 -56 73201
rect 56 74177 102 74189
rect 56 73201 62 74177
rect 96 73201 102 74177
rect 56 73189 102 73201
rect -46 73151 46 73157
rect -46 73117 -34 73151
rect 34 73117 46 73151
rect -46 73111 46 73117
rect -46 73043 46 73049
rect -46 73009 -34 73043
rect 34 73009 46 73043
rect -46 73003 46 73009
rect -102 72959 -56 72971
rect -102 71983 -96 72959
rect -62 71983 -56 72959
rect -102 71971 -56 71983
rect 56 72959 102 72971
rect 56 71983 62 72959
rect 96 71983 102 72959
rect 56 71971 102 71983
rect -46 71933 46 71939
rect -46 71899 -34 71933
rect 34 71899 46 71933
rect -46 71893 46 71899
rect -46 71825 46 71831
rect -46 71791 -34 71825
rect 34 71791 46 71825
rect -46 71785 46 71791
rect -102 71741 -56 71753
rect -102 70765 -96 71741
rect -62 70765 -56 71741
rect -102 70753 -56 70765
rect 56 71741 102 71753
rect 56 70765 62 71741
rect 96 70765 102 71741
rect 56 70753 102 70765
rect -46 70715 46 70721
rect -46 70681 -34 70715
rect 34 70681 46 70715
rect -46 70675 46 70681
rect -46 70607 46 70613
rect -46 70573 -34 70607
rect 34 70573 46 70607
rect -46 70567 46 70573
rect -102 70523 -56 70535
rect -102 69547 -96 70523
rect -62 69547 -56 70523
rect -102 69535 -56 69547
rect 56 70523 102 70535
rect 56 69547 62 70523
rect 96 69547 102 70523
rect 56 69535 102 69547
rect -46 69497 46 69503
rect -46 69463 -34 69497
rect 34 69463 46 69497
rect -46 69457 46 69463
rect -46 69389 46 69395
rect -46 69355 -34 69389
rect 34 69355 46 69389
rect -46 69349 46 69355
rect -102 69305 -56 69317
rect -102 68329 -96 69305
rect -62 68329 -56 69305
rect -102 68317 -56 68329
rect 56 69305 102 69317
rect 56 68329 62 69305
rect 96 68329 102 69305
rect 56 68317 102 68329
rect -46 68279 46 68285
rect -46 68245 -34 68279
rect 34 68245 46 68279
rect -46 68239 46 68245
rect -46 68171 46 68177
rect -46 68137 -34 68171
rect 34 68137 46 68171
rect -46 68131 46 68137
rect -102 68087 -56 68099
rect -102 67111 -96 68087
rect -62 67111 -56 68087
rect -102 67099 -56 67111
rect 56 68087 102 68099
rect 56 67111 62 68087
rect 96 67111 102 68087
rect 56 67099 102 67111
rect -46 67061 46 67067
rect -46 67027 -34 67061
rect 34 67027 46 67061
rect -46 67021 46 67027
rect -46 66953 46 66959
rect -46 66919 -34 66953
rect 34 66919 46 66953
rect -46 66913 46 66919
rect -102 66869 -56 66881
rect -102 65893 -96 66869
rect -62 65893 -56 66869
rect -102 65881 -56 65893
rect 56 66869 102 66881
rect 56 65893 62 66869
rect 96 65893 102 66869
rect 56 65881 102 65893
rect -46 65843 46 65849
rect -46 65809 -34 65843
rect 34 65809 46 65843
rect -46 65803 46 65809
rect -46 65735 46 65741
rect -46 65701 -34 65735
rect 34 65701 46 65735
rect -46 65695 46 65701
rect -102 65651 -56 65663
rect -102 64675 -96 65651
rect -62 64675 -56 65651
rect -102 64663 -56 64675
rect 56 65651 102 65663
rect 56 64675 62 65651
rect 96 64675 102 65651
rect 56 64663 102 64675
rect -46 64625 46 64631
rect -46 64591 -34 64625
rect 34 64591 46 64625
rect -46 64585 46 64591
rect -46 64517 46 64523
rect -46 64483 -34 64517
rect 34 64483 46 64517
rect -46 64477 46 64483
rect -102 64433 -56 64445
rect -102 63457 -96 64433
rect -62 63457 -56 64433
rect -102 63445 -56 63457
rect 56 64433 102 64445
rect 56 63457 62 64433
rect 96 63457 102 64433
rect 56 63445 102 63457
rect -46 63407 46 63413
rect -46 63373 -34 63407
rect 34 63373 46 63407
rect -46 63367 46 63373
rect -46 63299 46 63305
rect -46 63265 -34 63299
rect 34 63265 46 63299
rect -46 63259 46 63265
rect -102 63215 -56 63227
rect -102 62239 -96 63215
rect -62 62239 -56 63215
rect -102 62227 -56 62239
rect 56 63215 102 63227
rect 56 62239 62 63215
rect 96 62239 102 63215
rect 56 62227 102 62239
rect -46 62189 46 62195
rect -46 62155 -34 62189
rect 34 62155 46 62189
rect -46 62149 46 62155
rect -46 62081 46 62087
rect -46 62047 -34 62081
rect 34 62047 46 62081
rect -46 62041 46 62047
rect -102 61997 -56 62009
rect -102 61021 -96 61997
rect -62 61021 -56 61997
rect -102 61009 -56 61021
rect 56 61997 102 62009
rect 56 61021 62 61997
rect 96 61021 102 61997
rect 56 61009 102 61021
rect -46 60971 46 60977
rect -46 60937 -34 60971
rect 34 60937 46 60971
rect -46 60931 46 60937
rect -46 60863 46 60869
rect -46 60829 -34 60863
rect 34 60829 46 60863
rect -46 60823 46 60829
rect -102 60779 -56 60791
rect -102 59803 -96 60779
rect -62 59803 -56 60779
rect -102 59791 -56 59803
rect 56 60779 102 60791
rect 56 59803 62 60779
rect 96 59803 102 60779
rect 56 59791 102 59803
rect -46 59753 46 59759
rect -46 59719 -34 59753
rect 34 59719 46 59753
rect -46 59713 46 59719
rect -46 59645 46 59651
rect -46 59611 -34 59645
rect 34 59611 46 59645
rect -46 59605 46 59611
rect -102 59561 -56 59573
rect -102 58585 -96 59561
rect -62 58585 -56 59561
rect -102 58573 -56 58585
rect 56 59561 102 59573
rect 56 58585 62 59561
rect 96 58585 102 59561
rect 56 58573 102 58585
rect -46 58535 46 58541
rect -46 58501 -34 58535
rect 34 58501 46 58535
rect -46 58495 46 58501
rect -46 58427 46 58433
rect -46 58393 -34 58427
rect 34 58393 46 58427
rect -46 58387 46 58393
rect -102 58343 -56 58355
rect -102 57367 -96 58343
rect -62 57367 -56 58343
rect -102 57355 -56 57367
rect 56 58343 102 58355
rect 56 57367 62 58343
rect 96 57367 102 58343
rect 56 57355 102 57367
rect -46 57317 46 57323
rect -46 57283 -34 57317
rect 34 57283 46 57317
rect -46 57277 46 57283
rect -46 57209 46 57215
rect -46 57175 -34 57209
rect 34 57175 46 57209
rect -46 57169 46 57175
rect -102 57125 -56 57137
rect -102 56149 -96 57125
rect -62 56149 -56 57125
rect -102 56137 -56 56149
rect 56 57125 102 57137
rect 56 56149 62 57125
rect 96 56149 102 57125
rect 56 56137 102 56149
rect -46 56099 46 56105
rect -46 56065 -34 56099
rect 34 56065 46 56099
rect -46 56059 46 56065
rect -46 55991 46 55997
rect -46 55957 -34 55991
rect 34 55957 46 55991
rect -46 55951 46 55957
rect -102 55907 -56 55919
rect -102 54931 -96 55907
rect -62 54931 -56 55907
rect -102 54919 -56 54931
rect 56 55907 102 55919
rect 56 54931 62 55907
rect 96 54931 102 55907
rect 56 54919 102 54931
rect -46 54881 46 54887
rect -46 54847 -34 54881
rect 34 54847 46 54881
rect -46 54841 46 54847
rect -46 54773 46 54779
rect -46 54739 -34 54773
rect 34 54739 46 54773
rect -46 54733 46 54739
rect -102 54689 -56 54701
rect -102 53713 -96 54689
rect -62 53713 -56 54689
rect -102 53701 -56 53713
rect 56 54689 102 54701
rect 56 53713 62 54689
rect 96 53713 102 54689
rect 56 53701 102 53713
rect -46 53663 46 53669
rect -46 53629 -34 53663
rect 34 53629 46 53663
rect -46 53623 46 53629
rect -46 53555 46 53561
rect -46 53521 -34 53555
rect 34 53521 46 53555
rect -46 53515 46 53521
rect -102 53471 -56 53483
rect -102 52495 -96 53471
rect -62 52495 -56 53471
rect -102 52483 -56 52495
rect 56 53471 102 53483
rect 56 52495 62 53471
rect 96 52495 102 53471
rect 56 52483 102 52495
rect -46 52445 46 52451
rect -46 52411 -34 52445
rect 34 52411 46 52445
rect -46 52405 46 52411
rect -46 52337 46 52343
rect -46 52303 -34 52337
rect 34 52303 46 52337
rect -46 52297 46 52303
rect -102 52253 -56 52265
rect -102 51277 -96 52253
rect -62 51277 -56 52253
rect -102 51265 -56 51277
rect 56 52253 102 52265
rect 56 51277 62 52253
rect 96 51277 102 52253
rect 56 51265 102 51277
rect -46 51227 46 51233
rect -46 51193 -34 51227
rect 34 51193 46 51227
rect -46 51187 46 51193
rect -46 51119 46 51125
rect -46 51085 -34 51119
rect 34 51085 46 51119
rect -46 51079 46 51085
rect -102 51035 -56 51047
rect -102 50059 -96 51035
rect -62 50059 -56 51035
rect -102 50047 -56 50059
rect 56 51035 102 51047
rect 56 50059 62 51035
rect 96 50059 102 51035
rect 56 50047 102 50059
rect -46 50009 46 50015
rect -46 49975 -34 50009
rect 34 49975 46 50009
rect -46 49969 46 49975
rect -46 49901 46 49907
rect -46 49867 -34 49901
rect 34 49867 46 49901
rect -46 49861 46 49867
rect -102 49817 -56 49829
rect -102 48841 -96 49817
rect -62 48841 -56 49817
rect -102 48829 -56 48841
rect 56 49817 102 49829
rect 56 48841 62 49817
rect 96 48841 102 49817
rect 56 48829 102 48841
rect -46 48791 46 48797
rect -46 48757 -34 48791
rect 34 48757 46 48791
rect -46 48751 46 48757
rect -46 48683 46 48689
rect -46 48649 -34 48683
rect 34 48649 46 48683
rect -46 48643 46 48649
rect -102 48599 -56 48611
rect -102 47623 -96 48599
rect -62 47623 -56 48599
rect -102 47611 -56 47623
rect 56 48599 102 48611
rect 56 47623 62 48599
rect 96 47623 102 48599
rect 56 47611 102 47623
rect -46 47573 46 47579
rect -46 47539 -34 47573
rect 34 47539 46 47573
rect -46 47533 46 47539
rect -46 47465 46 47471
rect -46 47431 -34 47465
rect 34 47431 46 47465
rect -46 47425 46 47431
rect -102 47381 -56 47393
rect -102 46405 -96 47381
rect -62 46405 -56 47381
rect -102 46393 -56 46405
rect 56 47381 102 47393
rect 56 46405 62 47381
rect 96 46405 102 47381
rect 56 46393 102 46405
rect -46 46355 46 46361
rect -46 46321 -34 46355
rect 34 46321 46 46355
rect -46 46315 46 46321
rect -46 46247 46 46253
rect -46 46213 -34 46247
rect 34 46213 46 46247
rect -46 46207 46 46213
rect -102 46163 -56 46175
rect -102 45187 -96 46163
rect -62 45187 -56 46163
rect -102 45175 -56 45187
rect 56 46163 102 46175
rect 56 45187 62 46163
rect 96 45187 102 46163
rect 56 45175 102 45187
rect -46 45137 46 45143
rect -46 45103 -34 45137
rect 34 45103 46 45137
rect -46 45097 46 45103
rect -46 45029 46 45035
rect -46 44995 -34 45029
rect 34 44995 46 45029
rect -46 44989 46 44995
rect -102 44945 -56 44957
rect -102 43969 -96 44945
rect -62 43969 -56 44945
rect -102 43957 -56 43969
rect 56 44945 102 44957
rect 56 43969 62 44945
rect 96 43969 102 44945
rect 56 43957 102 43969
rect -46 43919 46 43925
rect -46 43885 -34 43919
rect 34 43885 46 43919
rect -46 43879 46 43885
rect -46 43811 46 43817
rect -46 43777 -34 43811
rect 34 43777 46 43811
rect -46 43771 46 43777
rect -102 43727 -56 43739
rect -102 42751 -96 43727
rect -62 42751 -56 43727
rect -102 42739 -56 42751
rect 56 43727 102 43739
rect 56 42751 62 43727
rect 96 42751 102 43727
rect 56 42739 102 42751
rect -46 42701 46 42707
rect -46 42667 -34 42701
rect 34 42667 46 42701
rect -46 42661 46 42667
rect -46 42593 46 42599
rect -46 42559 -34 42593
rect 34 42559 46 42593
rect -46 42553 46 42559
rect -102 42509 -56 42521
rect -102 41533 -96 42509
rect -62 41533 -56 42509
rect -102 41521 -56 41533
rect 56 42509 102 42521
rect 56 41533 62 42509
rect 96 41533 102 42509
rect 56 41521 102 41533
rect -46 41483 46 41489
rect -46 41449 -34 41483
rect 34 41449 46 41483
rect -46 41443 46 41449
rect -46 41375 46 41381
rect -46 41341 -34 41375
rect 34 41341 46 41375
rect -46 41335 46 41341
rect -102 41291 -56 41303
rect -102 40315 -96 41291
rect -62 40315 -56 41291
rect -102 40303 -56 40315
rect 56 41291 102 41303
rect 56 40315 62 41291
rect 96 40315 102 41291
rect 56 40303 102 40315
rect -46 40265 46 40271
rect -46 40231 -34 40265
rect 34 40231 46 40265
rect -46 40225 46 40231
rect -46 40157 46 40163
rect -46 40123 -34 40157
rect 34 40123 46 40157
rect -46 40117 46 40123
rect -102 40073 -56 40085
rect -102 39097 -96 40073
rect -62 39097 -56 40073
rect -102 39085 -56 39097
rect 56 40073 102 40085
rect 56 39097 62 40073
rect 96 39097 102 40073
rect 56 39085 102 39097
rect -46 39047 46 39053
rect -46 39013 -34 39047
rect 34 39013 46 39047
rect -46 39007 46 39013
rect -46 38939 46 38945
rect -46 38905 -34 38939
rect 34 38905 46 38939
rect -46 38899 46 38905
rect -102 38855 -56 38867
rect -102 37879 -96 38855
rect -62 37879 -56 38855
rect -102 37867 -56 37879
rect 56 38855 102 38867
rect 56 37879 62 38855
rect 96 37879 102 38855
rect 56 37867 102 37879
rect -46 37829 46 37835
rect -46 37795 -34 37829
rect 34 37795 46 37829
rect -46 37789 46 37795
rect -46 37721 46 37727
rect -46 37687 -34 37721
rect 34 37687 46 37721
rect -46 37681 46 37687
rect -102 37637 -56 37649
rect -102 36661 -96 37637
rect -62 36661 -56 37637
rect -102 36649 -56 36661
rect 56 37637 102 37649
rect 56 36661 62 37637
rect 96 36661 102 37637
rect 56 36649 102 36661
rect -46 36611 46 36617
rect -46 36577 -34 36611
rect 34 36577 46 36611
rect -46 36571 46 36577
rect -46 36503 46 36509
rect -46 36469 -34 36503
rect 34 36469 46 36503
rect -46 36463 46 36469
rect -102 36419 -56 36431
rect -102 35443 -96 36419
rect -62 35443 -56 36419
rect -102 35431 -56 35443
rect 56 36419 102 36431
rect 56 35443 62 36419
rect 96 35443 102 36419
rect 56 35431 102 35443
rect -46 35393 46 35399
rect -46 35359 -34 35393
rect 34 35359 46 35393
rect -46 35353 46 35359
rect -46 35285 46 35291
rect -46 35251 -34 35285
rect 34 35251 46 35285
rect -46 35245 46 35251
rect -102 35201 -56 35213
rect -102 34225 -96 35201
rect -62 34225 -56 35201
rect -102 34213 -56 34225
rect 56 35201 102 35213
rect 56 34225 62 35201
rect 96 34225 102 35201
rect 56 34213 102 34225
rect -46 34175 46 34181
rect -46 34141 -34 34175
rect 34 34141 46 34175
rect -46 34135 46 34141
rect -46 34067 46 34073
rect -46 34033 -34 34067
rect 34 34033 46 34067
rect -46 34027 46 34033
rect -102 33983 -56 33995
rect -102 33007 -96 33983
rect -62 33007 -56 33983
rect -102 32995 -56 33007
rect 56 33983 102 33995
rect 56 33007 62 33983
rect 96 33007 102 33983
rect 56 32995 102 33007
rect -46 32957 46 32963
rect -46 32923 -34 32957
rect 34 32923 46 32957
rect -46 32917 46 32923
rect -46 32849 46 32855
rect -46 32815 -34 32849
rect 34 32815 46 32849
rect -46 32809 46 32815
rect -102 32765 -56 32777
rect -102 31789 -96 32765
rect -62 31789 -56 32765
rect -102 31777 -56 31789
rect 56 32765 102 32777
rect 56 31789 62 32765
rect 96 31789 102 32765
rect 56 31777 102 31789
rect -46 31739 46 31745
rect -46 31705 -34 31739
rect 34 31705 46 31739
rect -46 31699 46 31705
rect -46 31631 46 31637
rect -46 31597 -34 31631
rect 34 31597 46 31631
rect -46 31591 46 31597
rect -102 31547 -56 31559
rect -102 30571 -96 31547
rect -62 30571 -56 31547
rect -102 30559 -56 30571
rect 56 31547 102 31559
rect 56 30571 62 31547
rect 96 30571 102 31547
rect 56 30559 102 30571
rect -46 30521 46 30527
rect -46 30487 -34 30521
rect 34 30487 46 30521
rect -46 30481 46 30487
rect -46 30413 46 30419
rect -46 30379 -34 30413
rect 34 30379 46 30413
rect -46 30373 46 30379
rect -102 30329 -56 30341
rect -102 29353 -96 30329
rect -62 29353 -56 30329
rect -102 29341 -56 29353
rect 56 30329 102 30341
rect 56 29353 62 30329
rect 96 29353 102 30329
rect 56 29341 102 29353
rect -46 29303 46 29309
rect -46 29269 -34 29303
rect 34 29269 46 29303
rect -46 29263 46 29269
rect -46 29195 46 29201
rect -46 29161 -34 29195
rect 34 29161 46 29195
rect -46 29155 46 29161
rect -102 29111 -56 29123
rect -102 28135 -96 29111
rect -62 28135 -56 29111
rect -102 28123 -56 28135
rect 56 29111 102 29123
rect 56 28135 62 29111
rect 96 28135 102 29111
rect 56 28123 102 28135
rect -46 28085 46 28091
rect -46 28051 -34 28085
rect 34 28051 46 28085
rect -46 28045 46 28051
rect -46 27977 46 27983
rect -46 27943 -34 27977
rect 34 27943 46 27977
rect -46 27937 46 27943
rect -102 27893 -56 27905
rect -102 26917 -96 27893
rect -62 26917 -56 27893
rect -102 26905 -56 26917
rect 56 27893 102 27905
rect 56 26917 62 27893
rect 96 26917 102 27893
rect 56 26905 102 26917
rect -46 26867 46 26873
rect -46 26833 -34 26867
rect 34 26833 46 26867
rect -46 26827 46 26833
rect -46 26759 46 26765
rect -46 26725 -34 26759
rect 34 26725 46 26759
rect -46 26719 46 26725
rect -102 26675 -56 26687
rect -102 25699 -96 26675
rect -62 25699 -56 26675
rect -102 25687 -56 25699
rect 56 26675 102 26687
rect 56 25699 62 26675
rect 96 25699 102 26675
rect 56 25687 102 25699
rect -46 25649 46 25655
rect -46 25615 -34 25649
rect 34 25615 46 25649
rect -46 25609 46 25615
rect -46 25541 46 25547
rect -46 25507 -34 25541
rect 34 25507 46 25541
rect -46 25501 46 25507
rect -102 25457 -56 25469
rect -102 24481 -96 25457
rect -62 24481 -56 25457
rect -102 24469 -56 24481
rect 56 25457 102 25469
rect 56 24481 62 25457
rect 96 24481 102 25457
rect 56 24469 102 24481
rect -46 24431 46 24437
rect -46 24397 -34 24431
rect 34 24397 46 24431
rect -46 24391 46 24397
rect -46 24323 46 24329
rect -46 24289 -34 24323
rect 34 24289 46 24323
rect -46 24283 46 24289
rect -102 24239 -56 24251
rect -102 23263 -96 24239
rect -62 23263 -56 24239
rect -102 23251 -56 23263
rect 56 24239 102 24251
rect 56 23263 62 24239
rect 96 23263 102 24239
rect 56 23251 102 23263
rect -46 23213 46 23219
rect -46 23179 -34 23213
rect 34 23179 46 23213
rect -46 23173 46 23179
rect -46 23105 46 23111
rect -46 23071 -34 23105
rect 34 23071 46 23105
rect -46 23065 46 23071
rect -102 23021 -56 23033
rect -102 22045 -96 23021
rect -62 22045 -56 23021
rect -102 22033 -56 22045
rect 56 23021 102 23033
rect 56 22045 62 23021
rect 96 22045 102 23021
rect 56 22033 102 22045
rect -46 21995 46 22001
rect -46 21961 -34 21995
rect 34 21961 46 21995
rect -46 21955 46 21961
rect -46 21887 46 21893
rect -46 21853 -34 21887
rect 34 21853 46 21887
rect -46 21847 46 21853
rect -102 21803 -56 21815
rect -102 20827 -96 21803
rect -62 20827 -56 21803
rect -102 20815 -56 20827
rect 56 21803 102 21815
rect 56 20827 62 21803
rect 96 20827 102 21803
rect 56 20815 102 20827
rect -46 20777 46 20783
rect -46 20743 -34 20777
rect 34 20743 46 20777
rect -46 20737 46 20743
rect -46 20669 46 20675
rect -46 20635 -34 20669
rect 34 20635 46 20669
rect -46 20629 46 20635
rect -102 20585 -56 20597
rect -102 19609 -96 20585
rect -62 19609 -56 20585
rect -102 19597 -56 19609
rect 56 20585 102 20597
rect 56 19609 62 20585
rect 96 19609 102 20585
rect 56 19597 102 19609
rect -46 19559 46 19565
rect -46 19525 -34 19559
rect 34 19525 46 19559
rect -46 19519 46 19525
rect -46 19451 46 19457
rect -46 19417 -34 19451
rect 34 19417 46 19451
rect -46 19411 46 19417
rect -102 19367 -56 19379
rect -102 18391 -96 19367
rect -62 18391 -56 19367
rect -102 18379 -56 18391
rect 56 19367 102 19379
rect 56 18391 62 19367
rect 96 18391 102 19367
rect 56 18379 102 18391
rect -46 18341 46 18347
rect -46 18307 -34 18341
rect 34 18307 46 18341
rect -46 18301 46 18307
rect -46 18233 46 18239
rect -46 18199 -34 18233
rect 34 18199 46 18233
rect -46 18193 46 18199
rect -102 18149 -56 18161
rect -102 17173 -96 18149
rect -62 17173 -56 18149
rect -102 17161 -56 17173
rect 56 18149 102 18161
rect 56 17173 62 18149
rect 96 17173 102 18149
rect 56 17161 102 17173
rect -46 17123 46 17129
rect -46 17089 -34 17123
rect 34 17089 46 17123
rect -46 17083 46 17089
rect -46 17015 46 17021
rect -46 16981 -34 17015
rect 34 16981 46 17015
rect -46 16975 46 16981
rect -102 16931 -56 16943
rect -102 15955 -96 16931
rect -62 15955 -56 16931
rect -102 15943 -56 15955
rect 56 16931 102 16943
rect 56 15955 62 16931
rect 96 15955 102 16931
rect 56 15943 102 15955
rect -46 15905 46 15911
rect -46 15871 -34 15905
rect 34 15871 46 15905
rect -46 15865 46 15871
rect -46 15797 46 15803
rect -46 15763 -34 15797
rect 34 15763 46 15797
rect -46 15757 46 15763
rect -102 15713 -56 15725
rect -102 14737 -96 15713
rect -62 14737 -56 15713
rect -102 14725 -56 14737
rect 56 15713 102 15725
rect 56 14737 62 15713
rect 96 14737 102 15713
rect 56 14725 102 14737
rect -46 14687 46 14693
rect -46 14653 -34 14687
rect 34 14653 46 14687
rect -46 14647 46 14653
rect -46 14579 46 14585
rect -46 14545 -34 14579
rect 34 14545 46 14579
rect -46 14539 46 14545
rect -102 14495 -56 14507
rect -102 13519 -96 14495
rect -62 13519 -56 14495
rect -102 13507 -56 13519
rect 56 14495 102 14507
rect 56 13519 62 14495
rect 96 13519 102 14495
rect 56 13507 102 13519
rect -46 13469 46 13475
rect -46 13435 -34 13469
rect 34 13435 46 13469
rect -46 13429 46 13435
rect -46 13361 46 13367
rect -46 13327 -34 13361
rect 34 13327 46 13361
rect -46 13321 46 13327
rect -102 13277 -56 13289
rect -102 12301 -96 13277
rect -62 12301 -56 13277
rect -102 12289 -56 12301
rect 56 13277 102 13289
rect 56 12301 62 13277
rect 96 12301 102 13277
rect 56 12289 102 12301
rect -46 12251 46 12257
rect -46 12217 -34 12251
rect 34 12217 46 12251
rect -46 12211 46 12217
rect -46 12143 46 12149
rect -46 12109 -34 12143
rect 34 12109 46 12143
rect -46 12103 46 12109
rect -102 12059 -56 12071
rect -102 11083 -96 12059
rect -62 11083 -56 12059
rect -102 11071 -56 11083
rect 56 12059 102 12071
rect 56 11083 62 12059
rect 96 11083 102 12059
rect 56 11071 102 11083
rect -46 11033 46 11039
rect -46 10999 -34 11033
rect 34 10999 46 11033
rect -46 10993 46 10999
rect -46 10925 46 10931
rect -46 10891 -34 10925
rect 34 10891 46 10925
rect -46 10885 46 10891
rect -102 10841 -56 10853
rect -102 9865 -96 10841
rect -62 9865 -56 10841
rect -102 9853 -56 9865
rect 56 10841 102 10853
rect 56 9865 62 10841
rect 96 9865 102 10841
rect 56 9853 102 9865
rect -46 9815 46 9821
rect -46 9781 -34 9815
rect 34 9781 46 9815
rect -46 9775 46 9781
rect -46 9707 46 9713
rect -46 9673 -34 9707
rect 34 9673 46 9707
rect -46 9667 46 9673
rect -102 9623 -56 9635
rect -102 8647 -96 9623
rect -62 8647 -56 9623
rect -102 8635 -56 8647
rect 56 9623 102 9635
rect 56 8647 62 9623
rect 96 8647 102 9623
rect 56 8635 102 8647
rect -46 8597 46 8603
rect -46 8563 -34 8597
rect 34 8563 46 8597
rect -46 8557 46 8563
rect -46 8489 46 8495
rect -46 8455 -34 8489
rect 34 8455 46 8489
rect -46 8449 46 8455
rect -102 8405 -56 8417
rect -102 7429 -96 8405
rect -62 7429 -56 8405
rect -102 7417 -56 7429
rect 56 8405 102 8417
rect 56 7429 62 8405
rect 96 7429 102 8405
rect 56 7417 102 7429
rect -46 7379 46 7385
rect -46 7345 -34 7379
rect 34 7345 46 7379
rect -46 7339 46 7345
rect -46 7271 46 7277
rect -46 7237 -34 7271
rect 34 7237 46 7271
rect -46 7231 46 7237
rect -102 7187 -56 7199
rect -102 6211 -96 7187
rect -62 6211 -56 7187
rect -102 6199 -56 6211
rect 56 7187 102 7199
rect 56 6211 62 7187
rect 96 6211 102 7187
rect 56 6199 102 6211
rect -46 6161 46 6167
rect -46 6127 -34 6161
rect 34 6127 46 6161
rect -46 6121 46 6127
rect -46 6053 46 6059
rect -46 6019 -34 6053
rect 34 6019 46 6053
rect -46 6013 46 6019
rect -102 5969 -56 5981
rect -102 4993 -96 5969
rect -62 4993 -56 5969
rect -102 4981 -56 4993
rect 56 5969 102 5981
rect 56 4993 62 5969
rect 96 4993 102 5969
rect 56 4981 102 4993
rect -46 4943 46 4949
rect -46 4909 -34 4943
rect 34 4909 46 4943
rect -46 4903 46 4909
rect -46 4835 46 4841
rect -46 4801 -34 4835
rect 34 4801 46 4835
rect -46 4795 46 4801
rect -102 4751 -56 4763
rect -102 3775 -96 4751
rect -62 3775 -56 4751
rect -102 3763 -56 3775
rect 56 4751 102 4763
rect 56 3775 62 4751
rect 96 3775 102 4751
rect 56 3763 102 3775
rect -46 3725 46 3731
rect -46 3691 -34 3725
rect 34 3691 46 3725
rect -46 3685 46 3691
rect -46 3617 46 3623
rect -46 3583 -34 3617
rect 34 3583 46 3617
rect -46 3577 46 3583
rect -102 3533 -56 3545
rect -102 2557 -96 3533
rect -62 2557 -56 3533
rect -102 2545 -56 2557
rect 56 3533 102 3545
rect 56 2557 62 3533
rect 96 2557 102 3533
rect 56 2545 102 2557
rect -46 2507 46 2513
rect -46 2473 -34 2507
rect 34 2473 46 2507
rect -46 2467 46 2473
rect -46 2399 46 2405
rect -46 2365 -34 2399
rect 34 2365 46 2399
rect -46 2359 46 2365
rect -102 2315 -56 2327
rect -102 1339 -96 2315
rect -62 1339 -56 2315
rect -102 1327 -56 1339
rect 56 2315 102 2327
rect 56 1339 62 2315
rect 96 1339 102 2315
rect 56 1327 102 1339
rect -46 1289 46 1295
rect -46 1255 -34 1289
rect 34 1255 46 1289
rect -46 1249 46 1255
rect -46 1181 46 1187
rect -46 1147 -34 1181
rect 34 1147 46 1181
rect -46 1141 46 1147
rect -102 1097 -56 1109
rect -102 121 -96 1097
rect -62 121 -56 1097
rect -102 109 -56 121
rect 56 1097 102 1109
rect 56 121 62 1097
rect 96 121 102 1097
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -1097 -96 -121
rect -62 -1097 -56 -121
rect -102 -1109 -56 -1097
rect 56 -121 102 -109
rect 56 -1097 62 -121
rect 96 -1097 102 -121
rect 56 -1109 102 -1097
rect -46 -1147 46 -1141
rect -46 -1181 -34 -1147
rect 34 -1181 46 -1147
rect -46 -1187 46 -1181
rect -46 -1255 46 -1249
rect -46 -1289 -34 -1255
rect 34 -1289 46 -1255
rect -46 -1295 46 -1289
rect -102 -1339 -56 -1327
rect -102 -2315 -96 -1339
rect -62 -2315 -56 -1339
rect -102 -2327 -56 -2315
rect 56 -1339 102 -1327
rect 56 -2315 62 -1339
rect 96 -2315 102 -1339
rect 56 -2327 102 -2315
rect -46 -2365 46 -2359
rect -46 -2399 -34 -2365
rect 34 -2399 46 -2365
rect -46 -2405 46 -2399
rect -46 -2473 46 -2467
rect -46 -2507 -34 -2473
rect 34 -2507 46 -2473
rect -46 -2513 46 -2507
rect -102 -2557 -56 -2545
rect -102 -3533 -96 -2557
rect -62 -3533 -56 -2557
rect -102 -3545 -56 -3533
rect 56 -2557 102 -2545
rect 56 -3533 62 -2557
rect 96 -3533 102 -2557
rect 56 -3545 102 -3533
rect -46 -3583 46 -3577
rect -46 -3617 -34 -3583
rect 34 -3617 46 -3583
rect -46 -3623 46 -3617
rect -46 -3691 46 -3685
rect -46 -3725 -34 -3691
rect 34 -3725 46 -3691
rect -46 -3731 46 -3725
rect -102 -3775 -56 -3763
rect -102 -4751 -96 -3775
rect -62 -4751 -56 -3775
rect -102 -4763 -56 -4751
rect 56 -3775 102 -3763
rect 56 -4751 62 -3775
rect 96 -4751 102 -3775
rect 56 -4763 102 -4751
rect -46 -4801 46 -4795
rect -46 -4835 -34 -4801
rect 34 -4835 46 -4801
rect -46 -4841 46 -4835
rect -46 -4909 46 -4903
rect -46 -4943 -34 -4909
rect 34 -4943 46 -4909
rect -46 -4949 46 -4943
rect -102 -4993 -56 -4981
rect -102 -5969 -96 -4993
rect -62 -5969 -56 -4993
rect -102 -5981 -56 -5969
rect 56 -4993 102 -4981
rect 56 -5969 62 -4993
rect 96 -5969 102 -4993
rect 56 -5981 102 -5969
rect -46 -6019 46 -6013
rect -46 -6053 -34 -6019
rect 34 -6053 46 -6019
rect -46 -6059 46 -6053
rect -46 -6127 46 -6121
rect -46 -6161 -34 -6127
rect 34 -6161 46 -6127
rect -46 -6167 46 -6161
rect -102 -6211 -56 -6199
rect -102 -7187 -96 -6211
rect -62 -7187 -56 -6211
rect -102 -7199 -56 -7187
rect 56 -6211 102 -6199
rect 56 -7187 62 -6211
rect 96 -7187 102 -6211
rect 56 -7199 102 -7187
rect -46 -7237 46 -7231
rect -46 -7271 -34 -7237
rect 34 -7271 46 -7237
rect -46 -7277 46 -7271
rect -46 -7345 46 -7339
rect -46 -7379 -34 -7345
rect 34 -7379 46 -7345
rect -46 -7385 46 -7379
rect -102 -7429 -56 -7417
rect -102 -8405 -96 -7429
rect -62 -8405 -56 -7429
rect -102 -8417 -56 -8405
rect 56 -7429 102 -7417
rect 56 -8405 62 -7429
rect 96 -8405 102 -7429
rect 56 -8417 102 -8405
rect -46 -8455 46 -8449
rect -46 -8489 -34 -8455
rect 34 -8489 46 -8455
rect -46 -8495 46 -8489
rect -46 -8563 46 -8557
rect -46 -8597 -34 -8563
rect 34 -8597 46 -8563
rect -46 -8603 46 -8597
rect -102 -8647 -56 -8635
rect -102 -9623 -96 -8647
rect -62 -9623 -56 -8647
rect -102 -9635 -56 -9623
rect 56 -8647 102 -8635
rect 56 -9623 62 -8647
rect 96 -9623 102 -8647
rect 56 -9635 102 -9623
rect -46 -9673 46 -9667
rect -46 -9707 -34 -9673
rect 34 -9707 46 -9673
rect -46 -9713 46 -9707
rect -46 -9781 46 -9775
rect -46 -9815 -34 -9781
rect 34 -9815 46 -9781
rect -46 -9821 46 -9815
rect -102 -9865 -56 -9853
rect -102 -10841 -96 -9865
rect -62 -10841 -56 -9865
rect -102 -10853 -56 -10841
rect 56 -9865 102 -9853
rect 56 -10841 62 -9865
rect 96 -10841 102 -9865
rect 56 -10853 102 -10841
rect -46 -10891 46 -10885
rect -46 -10925 -34 -10891
rect 34 -10925 46 -10891
rect -46 -10931 46 -10925
rect -46 -10999 46 -10993
rect -46 -11033 -34 -10999
rect 34 -11033 46 -10999
rect -46 -11039 46 -11033
rect -102 -11083 -56 -11071
rect -102 -12059 -96 -11083
rect -62 -12059 -56 -11083
rect -102 -12071 -56 -12059
rect 56 -11083 102 -11071
rect 56 -12059 62 -11083
rect 96 -12059 102 -11083
rect 56 -12071 102 -12059
rect -46 -12109 46 -12103
rect -46 -12143 -34 -12109
rect 34 -12143 46 -12109
rect -46 -12149 46 -12143
rect -46 -12217 46 -12211
rect -46 -12251 -34 -12217
rect 34 -12251 46 -12217
rect -46 -12257 46 -12251
rect -102 -12301 -56 -12289
rect -102 -13277 -96 -12301
rect -62 -13277 -56 -12301
rect -102 -13289 -56 -13277
rect 56 -12301 102 -12289
rect 56 -13277 62 -12301
rect 96 -13277 102 -12301
rect 56 -13289 102 -13277
rect -46 -13327 46 -13321
rect -46 -13361 -34 -13327
rect 34 -13361 46 -13327
rect -46 -13367 46 -13361
rect -46 -13435 46 -13429
rect -46 -13469 -34 -13435
rect 34 -13469 46 -13435
rect -46 -13475 46 -13469
rect -102 -13519 -56 -13507
rect -102 -14495 -96 -13519
rect -62 -14495 -56 -13519
rect -102 -14507 -56 -14495
rect 56 -13519 102 -13507
rect 56 -14495 62 -13519
rect 96 -14495 102 -13519
rect 56 -14507 102 -14495
rect -46 -14545 46 -14539
rect -46 -14579 -34 -14545
rect 34 -14579 46 -14545
rect -46 -14585 46 -14579
rect -46 -14653 46 -14647
rect -46 -14687 -34 -14653
rect 34 -14687 46 -14653
rect -46 -14693 46 -14687
rect -102 -14737 -56 -14725
rect -102 -15713 -96 -14737
rect -62 -15713 -56 -14737
rect -102 -15725 -56 -15713
rect 56 -14737 102 -14725
rect 56 -15713 62 -14737
rect 96 -15713 102 -14737
rect 56 -15725 102 -15713
rect -46 -15763 46 -15757
rect -46 -15797 -34 -15763
rect 34 -15797 46 -15763
rect -46 -15803 46 -15797
rect -46 -15871 46 -15865
rect -46 -15905 -34 -15871
rect 34 -15905 46 -15871
rect -46 -15911 46 -15905
rect -102 -15955 -56 -15943
rect -102 -16931 -96 -15955
rect -62 -16931 -56 -15955
rect -102 -16943 -56 -16931
rect 56 -15955 102 -15943
rect 56 -16931 62 -15955
rect 96 -16931 102 -15955
rect 56 -16943 102 -16931
rect -46 -16981 46 -16975
rect -46 -17015 -34 -16981
rect 34 -17015 46 -16981
rect -46 -17021 46 -17015
rect -46 -17089 46 -17083
rect -46 -17123 -34 -17089
rect 34 -17123 46 -17089
rect -46 -17129 46 -17123
rect -102 -17173 -56 -17161
rect -102 -18149 -96 -17173
rect -62 -18149 -56 -17173
rect -102 -18161 -56 -18149
rect 56 -17173 102 -17161
rect 56 -18149 62 -17173
rect 96 -18149 102 -17173
rect 56 -18161 102 -18149
rect -46 -18199 46 -18193
rect -46 -18233 -34 -18199
rect 34 -18233 46 -18199
rect -46 -18239 46 -18233
rect -46 -18307 46 -18301
rect -46 -18341 -34 -18307
rect 34 -18341 46 -18307
rect -46 -18347 46 -18341
rect -102 -18391 -56 -18379
rect -102 -19367 -96 -18391
rect -62 -19367 -56 -18391
rect -102 -19379 -56 -19367
rect 56 -18391 102 -18379
rect 56 -19367 62 -18391
rect 96 -19367 102 -18391
rect 56 -19379 102 -19367
rect -46 -19417 46 -19411
rect -46 -19451 -34 -19417
rect 34 -19451 46 -19417
rect -46 -19457 46 -19451
rect -46 -19525 46 -19519
rect -46 -19559 -34 -19525
rect 34 -19559 46 -19525
rect -46 -19565 46 -19559
rect -102 -19609 -56 -19597
rect -102 -20585 -96 -19609
rect -62 -20585 -56 -19609
rect -102 -20597 -56 -20585
rect 56 -19609 102 -19597
rect 56 -20585 62 -19609
rect 96 -20585 102 -19609
rect 56 -20597 102 -20585
rect -46 -20635 46 -20629
rect -46 -20669 -34 -20635
rect 34 -20669 46 -20635
rect -46 -20675 46 -20669
rect -46 -20743 46 -20737
rect -46 -20777 -34 -20743
rect 34 -20777 46 -20743
rect -46 -20783 46 -20777
rect -102 -20827 -56 -20815
rect -102 -21803 -96 -20827
rect -62 -21803 -56 -20827
rect -102 -21815 -56 -21803
rect 56 -20827 102 -20815
rect 56 -21803 62 -20827
rect 96 -21803 102 -20827
rect 56 -21815 102 -21803
rect -46 -21853 46 -21847
rect -46 -21887 -34 -21853
rect 34 -21887 46 -21853
rect -46 -21893 46 -21887
rect -46 -21961 46 -21955
rect -46 -21995 -34 -21961
rect 34 -21995 46 -21961
rect -46 -22001 46 -21995
rect -102 -22045 -56 -22033
rect -102 -23021 -96 -22045
rect -62 -23021 -56 -22045
rect -102 -23033 -56 -23021
rect 56 -22045 102 -22033
rect 56 -23021 62 -22045
rect 96 -23021 102 -22045
rect 56 -23033 102 -23021
rect -46 -23071 46 -23065
rect -46 -23105 -34 -23071
rect 34 -23105 46 -23071
rect -46 -23111 46 -23105
rect -46 -23179 46 -23173
rect -46 -23213 -34 -23179
rect 34 -23213 46 -23179
rect -46 -23219 46 -23213
rect -102 -23263 -56 -23251
rect -102 -24239 -96 -23263
rect -62 -24239 -56 -23263
rect -102 -24251 -56 -24239
rect 56 -23263 102 -23251
rect 56 -24239 62 -23263
rect 96 -24239 102 -23263
rect 56 -24251 102 -24239
rect -46 -24289 46 -24283
rect -46 -24323 -34 -24289
rect 34 -24323 46 -24289
rect -46 -24329 46 -24323
rect -46 -24397 46 -24391
rect -46 -24431 -34 -24397
rect 34 -24431 46 -24397
rect -46 -24437 46 -24431
rect -102 -24481 -56 -24469
rect -102 -25457 -96 -24481
rect -62 -25457 -56 -24481
rect -102 -25469 -56 -25457
rect 56 -24481 102 -24469
rect 56 -25457 62 -24481
rect 96 -25457 102 -24481
rect 56 -25469 102 -25457
rect -46 -25507 46 -25501
rect -46 -25541 -34 -25507
rect 34 -25541 46 -25507
rect -46 -25547 46 -25541
rect -46 -25615 46 -25609
rect -46 -25649 -34 -25615
rect 34 -25649 46 -25615
rect -46 -25655 46 -25649
rect -102 -25699 -56 -25687
rect -102 -26675 -96 -25699
rect -62 -26675 -56 -25699
rect -102 -26687 -56 -26675
rect 56 -25699 102 -25687
rect 56 -26675 62 -25699
rect 96 -26675 102 -25699
rect 56 -26687 102 -26675
rect -46 -26725 46 -26719
rect -46 -26759 -34 -26725
rect 34 -26759 46 -26725
rect -46 -26765 46 -26759
rect -46 -26833 46 -26827
rect -46 -26867 -34 -26833
rect 34 -26867 46 -26833
rect -46 -26873 46 -26867
rect -102 -26917 -56 -26905
rect -102 -27893 -96 -26917
rect -62 -27893 -56 -26917
rect -102 -27905 -56 -27893
rect 56 -26917 102 -26905
rect 56 -27893 62 -26917
rect 96 -27893 102 -26917
rect 56 -27905 102 -27893
rect -46 -27943 46 -27937
rect -46 -27977 -34 -27943
rect 34 -27977 46 -27943
rect -46 -27983 46 -27977
rect -46 -28051 46 -28045
rect -46 -28085 -34 -28051
rect 34 -28085 46 -28051
rect -46 -28091 46 -28085
rect -102 -28135 -56 -28123
rect -102 -29111 -96 -28135
rect -62 -29111 -56 -28135
rect -102 -29123 -56 -29111
rect 56 -28135 102 -28123
rect 56 -29111 62 -28135
rect 96 -29111 102 -28135
rect 56 -29123 102 -29111
rect -46 -29161 46 -29155
rect -46 -29195 -34 -29161
rect 34 -29195 46 -29161
rect -46 -29201 46 -29195
rect -46 -29269 46 -29263
rect -46 -29303 -34 -29269
rect 34 -29303 46 -29269
rect -46 -29309 46 -29303
rect -102 -29353 -56 -29341
rect -102 -30329 -96 -29353
rect -62 -30329 -56 -29353
rect -102 -30341 -56 -30329
rect 56 -29353 102 -29341
rect 56 -30329 62 -29353
rect 96 -30329 102 -29353
rect 56 -30341 102 -30329
rect -46 -30379 46 -30373
rect -46 -30413 -34 -30379
rect 34 -30413 46 -30379
rect -46 -30419 46 -30413
rect -46 -30487 46 -30481
rect -46 -30521 -34 -30487
rect 34 -30521 46 -30487
rect -46 -30527 46 -30521
rect -102 -30571 -56 -30559
rect -102 -31547 -96 -30571
rect -62 -31547 -56 -30571
rect -102 -31559 -56 -31547
rect 56 -30571 102 -30559
rect 56 -31547 62 -30571
rect 96 -31547 102 -30571
rect 56 -31559 102 -31547
rect -46 -31597 46 -31591
rect -46 -31631 -34 -31597
rect 34 -31631 46 -31597
rect -46 -31637 46 -31631
rect -46 -31705 46 -31699
rect -46 -31739 -34 -31705
rect 34 -31739 46 -31705
rect -46 -31745 46 -31739
rect -102 -31789 -56 -31777
rect -102 -32765 -96 -31789
rect -62 -32765 -56 -31789
rect -102 -32777 -56 -32765
rect 56 -31789 102 -31777
rect 56 -32765 62 -31789
rect 96 -32765 102 -31789
rect 56 -32777 102 -32765
rect -46 -32815 46 -32809
rect -46 -32849 -34 -32815
rect 34 -32849 46 -32815
rect -46 -32855 46 -32849
rect -46 -32923 46 -32917
rect -46 -32957 -34 -32923
rect 34 -32957 46 -32923
rect -46 -32963 46 -32957
rect -102 -33007 -56 -32995
rect -102 -33983 -96 -33007
rect -62 -33983 -56 -33007
rect -102 -33995 -56 -33983
rect 56 -33007 102 -32995
rect 56 -33983 62 -33007
rect 96 -33983 102 -33007
rect 56 -33995 102 -33983
rect -46 -34033 46 -34027
rect -46 -34067 -34 -34033
rect 34 -34067 46 -34033
rect -46 -34073 46 -34067
rect -46 -34141 46 -34135
rect -46 -34175 -34 -34141
rect 34 -34175 46 -34141
rect -46 -34181 46 -34175
rect -102 -34225 -56 -34213
rect -102 -35201 -96 -34225
rect -62 -35201 -56 -34225
rect -102 -35213 -56 -35201
rect 56 -34225 102 -34213
rect 56 -35201 62 -34225
rect 96 -35201 102 -34225
rect 56 -35213 102 -35201
rect -46 -35251 46 -35245
rect -46 -35285 -34 -35251
rect 34 -35285 46 -35251
rect -46 -35291 46 -35285
rect -46 -35359 46 -35353
rect -46 -35393 -34 -35359
rect 34 -35393 46 -35359
rect -46 -35399 46 -35393
rect -102 -35443 -56 -35431
rect -102 -36419 -96 -35443
rect -62 -36419 -56 -35443
rect -102 -36431 -56 -36419
rect 56 -35443 102 -35431
rect 56 -36419 62 -35443
rect 96 -36419 102 -35443
rect 56 -36431 102 -36419
rect -46 -36469 46 -36463
rect -46 -36503 -34 -36469
rect 34 -36503 46 -36469
rect -46 -36509 46 -36503
rect -46 -36577 46 -36571
rect -46 -36611 -34 -36577
rect 34 -36611 46 -36577
rect -46 -36617 46 -36611
rect -102 -36661 -56 -36649
rect -102 -37637 -96 -36661
rect -62 -37637 -56 -36661
rect -102 -37649 -56 -37637
rect 56 -36661 102 -36649
rect 56 -37637 62 -36661
rect 96 -37637 102 -36661
rect 56 -37649 102 -37637
rect -46 -37687 46 -37681
rect -46 -37721 -34 -37687
rect 34 -37721 46 -37687
rect -46 -37727 46 -37721
rect -46 -37795 46 -37789
rect -46 -37829 -34 -37795
rect 34 -37829 46 -37795
rect -46 -37835 46 -37829
rect -102 -37879 -56 -37867
rect -102 -38855 -96 -37879
rect -62 -38855 -56 -37879
rect -102 -38867 -56 -38855
rect 56 -37879 102 -37867
rect 56 -38855 62 -37879
rect 96 -38855 102 -37879
rect 56 -38867 102 -38855
rect -46 -38905 46 -38899
rect -46 -38939 -34 -38905
rect 34 -38939 46 -38905
rect -46 -38945 46 -38939
rect -46 -39013 46 -39007
rect -46 -39047 -34 -39013
rect 34 -39047 46 -39013
rect -46 -39053 46 -39047
rect -102 -39097 -56 -39085
rect -102 -40073 -96 -39097
rect -62 -40073 -56 -39097
rect -102 -40085 -56 -40073
rect 56 -39097 102 -39085
rect 56 -40073 62 -39097
rect 96 -40073 102 -39097
rect 56 -40085 102 -40073
rect -46 -40123 46 -40117
rect -46 -40157 -34 -40123
rect 34 -40157 46 -40123
rect -46 -40163 46 -40157
rect -46 -40231 46 -40225
rect -46 -40265 -34 -40231
rect 34 -40265 46 -40231
rect -46 -40271 46 -40265
rect -102 -40315 -56 -40303
rect -102 -41291 -96 -40315
rect -62 -41291 -56 -40315
rect -102 -41303 -56 -41291
rect 56 -40315 102 -40303
rect 56 -41291 62 -40315
rect 96 -41291 102 -40315
rect 56 -41303 102 -41291
rect -46 -41341 46 -41335
rect -46 -41375 -34 -41341
rect 34 -41375 46 -41341
rect -46 -41381 46 -41375
rect -46 -41449 46 -41443
rect -46 -41483 -34 -41449
rect 34 -41483 46 -41449
rect -46 -41489 46 -41483
rect -102 -41533 -56 -41521
rect -102 -42509 -96 -41533
rect -62 -42509 -56 -41533
rect -102 -42521 -56 -42509
rect 56 -41533 102 -41521
rect 56 -42509 62 -41533
rect 96 -42509 102 -41533
rect 56 -42521 102 -42509
rect -46 -42559 46 -42553
rect -46 -42593 -34 -42559
rect 34 -42593 46 -42559
rect -46 -42599 46 -42593
rect -46 -42667 46 -42661
rect -46 -42701 -34 -42667
rect 34 -42701 46 -42667
rect -46 -42707 46 -42701
rect -102 -42751 -56 -42739
rect -102 -43727 -96 -42751
rect -62 -43727 -56 -42751
rect -102 -43739 -56 -43727
rect 56 -42751 102 -42739
rect 56 -43727 62 -42751
rect 96 -43727 102 -42751
rect 56 -43739 102 -43727
rect -46 -43777 46 -43771
rect -46 -43811 -34 -43777
rect 34 -43811 46 -43777
rect -46 -43817 46 -43811
rect -46 -43885 46 -43879
rect -46 -43919 -34 -43885
rect 34 -43919 46 -43885
rect -46 -43925 46 -43919
rect -102 -43969 -56 -43957
rect -102 -44945 -96 -43969
rect -62 -44945 -56 -43969
rect -102 -44957 -56 -44945
rect 56 -43969 102 -43957
rect 56 -44945 62 -43969
rect 96 -44945 102 -43969
rect 56 -44957 102 -44945
rect -46 -44995 46 -44989
rect -46 -45029 -34 -44995
rect 34 -45029 46 -44995
rect -46 -45035 46 -45029
rect -46 -45103 46 -45097
rect -46 -45137 -34 -45103
rect 34 -45137 46 -45103
rect -46 -45143 46 -45137
rect -102 -45187 -56 -45175
rect -102 -46163 -96 -45187
rect -62 -46163 -56 -45187
rect -102 -46175 -56 -46163
rect 56 -45187 102 -45175
rect 56 -46163 62 -45187
rect 96 -46163 102 -45187
rect 56 -46175 102 -46163
rect -46 -46213 46 -46207
rect -46 -46247 -34 -46213
rect 34 -46247 46 -46213
rect -46 -46253 46 -46247
rect -46 -46321 46 -46315
rect -46 -46355 -34 -46321
rect 34 -46355 46 -46321
rect -46 -46361 46 -46355
rect -102 -46405 -56 -46393
rect -102 -47381 -96 -46405
rect -62 -47381 -56 -46405
rect -102 -47393 -56 -47381
rect 56 -46405 102 -46393
rect 56 -47381 62 -46405
rect 96 -47381 102 -46405
rect 56 -47393 102 -47381
rect -46 -47431 46 -47425
rect -46 -47465 -34 -47431
rect 34 -47465 46 -47431
rect -46 -47471 46 -47465
rect -46 -47539 46 -47533
rect -46 -47573 -34 -47539
rect 34 -47573 46 -47539
rect -46 -47579 46 -47573
rect -102 -47623 -56 -47611
rect -102 -48599 -96 -47623
rect -62 -48599 -56 -47623
rect -102 -48611 -56 -48599
rect 56 -47623 102 -47611
rect 56 -48599 62 -47623
rect 96 -48599 102 -47623
rect 56 -48611 102 -48599
rect -46 -48649 46 -48643
rect -46 -48683 -34 -48649
rect 34 -48683 46 -48649
rect -46 -48689 46 -48683
rect -46 -48757 46 -48751
rect -46 -48791 -34 -48757
rect 34 -48791 46 -48757
rect -46 -48797 46 -48791
rect -102 -48841 -56 -48829
rect -102 -49817 -96 -48841
rect -62 -49817 -56 -48841
rect -102 -49829 -56 -49817
rect 56 -48841 102 -48829
rect 56 -49817 62 -48841
rect 96 -49817 102 -48841
rect 56 -49829 102 -49817
rect -46 -49867 46 -49861
rect -46 -49901 -34 -49867
rect 34 -49901 46 -49867
rect -46 -49907 46 -49901
rect -46 -49975 46 -49969
rect -46 -50009 -34 -49975
rect 34 -50009 46 -49975
rect -46 -50015 46 -50009
rect -102 -50059 -56 -50047
rect -102 -51035 -96 -50059
rect -62 -51035 -56 -50059
rect -102 -51047 -56 -51035
rect 56 -50059 102 -50047
rect 56 -51035 62 -50059
rect 96 -51035 102 -50059
rect 56 -51047 102 -51035
rect -46 -51085 46 -51079
rect -46 -51119 -34 -51085
rect 34 -51119 46 -51085
rect -46 -51125 46 -51119
rect -46 -51193 46 -51187
rect -46 -51227 -34 -51193
rect 34 -51227 46 -51193
rect -46 -51233 46 -51227
rect -102 -51277 -56 -51265
rect -102 -52253 -96 -51277
rect -62 -52253 -56 -51277
rect -102 -52265 -56 -52253
rect 56 -51277 102 -51265
rect 56 -52253 62 -51277
rect 96 -52253 102 -51277
rect 56 -52265 102 -52253
rect -46 -52303 46 -52297
rect -46 -52337 -34 -52303
rect 34 -52337 46 -52303
rect -46 -52343 46 -52337
rect -46 -52411 46 -52405
rect -46 -52445 -34 -52411
rect 34 -52445 46 -52411
rect -46 -52451 46 -52445
rect -102 -52495 -56 -52483
rect -102 -53471 -96 -52495
rect -62 -53471 -56 -52495
rect -102 -53483 -56 -53471
rect 56 -52495 102 -52483
rect 56 -53471 62 -52495
rect 96 -53471 102 -52495
rect 56 -53483 102 -53471
rect -46 -53521 46 -53515
rect -46 -53555 -34 -53521
rect 34 -53555 46 -53521
rect -46 -53561 46 -53555
rect -46 -53629 46 -53623
rect -46 -53663 -34 -53629
rect 34 -53663 46 -53629
rect -46 -53669 46 -53663
rect -102 -53713 -56 -53701
rect -102 -54689 -96 -53713
rect -62 -54689 -56 -53713
rect -102 -54701 -56 -54689
rect 56 -53713 102 -53701
rect 56 -54689 62 -53713
rect 96 -54689 102 -53713
rect 56 -54701 102 -54689
rect -46 -54739 46 -54733
rect -46 -54773 -34 -54739
rect 34 -54773 46 -54739
rect -46 -54779 46 -54773
rect -46 -54847 46 -54841
rect -46 -54881 -34 -54847
rect 34 -54881 46 -54847
rect -46 -54887 46 -54881
rect -102 -54931 -56 -54919
rect -102 -55907 -96 -54931
rect -62 -55907 -56 -54931
rect -102 -55919 -56 -55907
rect 56 -54931 102 -54919
rect 56 -55907 62 -54931
rect 96 -55907 102 -54931
rect 56 -55919 102 -55907
rect -46 -55957 46 -55951
rect -46 -55991 -34 -55957
rect 34 -55991 46 -55957
rect -46 -55997 46 -55991
rect -46 -56065 46 -56059
rect -46 -56099 -34 -56065
rect 34 -56099 46 -56065
rect -46 -56105 46 -56099
rect -102 -56149 -56 -56137
rect -102 -57125 -96 -56149
rect -62 -57125 -56 -56149
rect -102 -57137 -56 -57125
rect 56 -56149 102 -56137
rect 56 -57125 62 -56149
rect 96 -57125 102 -56149
rect 56 -57137 102 -57125
rect -46 -57175 46 -57169
rect -46 -57209 -34 -57175
rect 34 -57209 46 -57175
rect -46 -57215 46 -57209
rect -46 -57283 46 -57277
rect -46 -57317 -34 -57283
rect 34 -57317 46 -57283
rect -46 -57323 46 -57317
rect -102 -57367 -56 -57355
rect -102 -58343 -96 -57367
rect -62 -58343 -56 -57367
rect -102 -58355 -56 -58343
rect 56 -57367 102 -57355
rect 56 -58343 62 -57367
rect 96 -58343 102 -57367
rect 56 -58355 102 -58343
rect -46 -58393 46 -58387
rect -46 -58427 -34 -58393
rect 34 -58427 46 -58393
rect -46 -58433 46 -58427
rect -46 -58501 46 -58495
rect -46 -58535 -34 -58501
rect 34 -58535 46 -58501
rect -46 -58541 46 -58535
rect -102 -58585 -56 -58573
rect -102 -59561 -96 -58585
rect -62 -59561 -56 -58585
rect -102 -59573 -56 -59561
rect 56 -58585 102 -58573
rect 56 -59561 62 -58585
rect 96 -59561 102 -58585
rect 56 -59573 102 -59561
rect -46 -59611 46 -59605
rect -46 -59645 -34 -59611
rect 34 -59645 46 -59611
rect -46 -59651 46 -59645
rect -46 -59719 46 -59713
rect -46 -59753 -34 -59719
rect 34 -59753 46 -59719
rect -46 -59759 46 -59753
rect -102 -59803 -56 -59791
rect -102 -60779 -96 -59803
rect -62 -60779 -56 -59803
rect -102 -60791 -56 -60779
rect 56 -59803 102 -59791
rect 56 -60779 62 -59803
rect 96 -60779 102 -59803
rect 56 -60791 102 -60779
rect -46 -60829 46 -60823
rect -46 -60863 -34 -60829
rect 34 -60863 46 -60829
rect -46 -60869 46 -60863
rect -46 -60937 46 -60931
rect -46 -60971 -34 -60937
rect 34 -60971 46 -60937
rect -46 -60977 46 -60971
rect -102 -61021 -56 -61009
rect -102 -61997 -96 -61021
rect -62 -61997 -56 -61021
rect -102 -62009 -56 -61997
rect 56 -61021 102 -61009
rect 56 -61997 62 -61021
rect 96 -61997 102 -61021
rect 56 -62009 102 -61997
rect -46 -62047 46 -62041
rect -46 -62081 -34 -62047
rect 34 -62081 46 -62047
rect -46 -62087 46 -62081
rect -46 -62155 46 -62149
rect -46 -62189 -34 -62155
rect 34 -62189 46 -62155
rect -46 -62195 46 -62189
rect -102 -62239 -56 -62227
rect -102 -63215 -96 -62239
rect -62 -63215 -56 -62239
rect -102 -63227 -56 -63215
rect 56 -62239 102 -62227
rect 56 -63215 62 -62239
rect 96 -63215 102 -62239
rect 56 -63227 102 -63215
rect -46 -63265 46 -63259
rect -46 -63299 -34 -63265
rect 34 -63299 46 -63265
rect -46 -63305 46 -63299
rect -46 -63373 46 -63367
rect -46 -63407 -34 -63373
rect 34 -63407 46 -63373
rect -46 -63413 46 -63407
rect -102 -63457 -56 -63445
rect -102 -64433 -96 -63457
rect -62 -64433 -56 -63457
rect -102 -64445 -56 -64433
rect 56 -63457 102 -63445
rect 56 -64433 62 -63457
rect 96 -64433 102 -63457
rect 56 -64445 102 -64433
rect -46 -64483 46 -64477
rect -46 -64517 -34 -64483
rect 34 -64517 46 -64483
rect -46 -64523 46 -64517
rect -46 -64591 46 -64585
rect -46 -64625 -34 -64591
rect 34 -64625 46 -64591
rect -46 -64631 46 -64625
rect -102 -64675 -56 -64663
rect -102 -65651 -96 -64675
rect -62 -65651 -56 -64675
rect -102 -65663 -56 -65651
rect 56 -64675 102 -64663
rect 56 -65651 62 -64675
rect 96 -65651 102 -64675
rect 56 -65663 102 -65651
rect -46 -65701 46 -65695
rect -46 -65735 -34 -65701
rect 34 -65735 46 -65701
rect -46 -65741 46 -65735
rect -46 -65809 46 -65803
rect -46 -65843 -34 -65809
rect 34 -65843 46 -65809
rect -46 -65849 46 -65843
rect -102 -65893 -56 -65881
rect -102 -66869 -96 -65893
rect -62 -66869 -56 -65893
rect -102 -66881 -56 -66869
rect 56 -65893 102 -65881
rect 56 -66869 62 -65893
rect 96 -66869 102 -65893
rect 56 -66881 102 -66869
rect -46 -66919 46 -66913
rect -46 -66953 -34 -66919
rect 34 -66953 46 -66919
rect -46 -66959 46 -66953
rect -46 -67027 46 -67021
rect -46 -67061 -34 -67027
rect 34 -67061 46 -67027
rect -46 -67067 46 -67061
rect -102 -67111 -56 -67099
rect -102 -68087 -96 -67111
rect -62 -68087 -56 -67111
rect -102 -68099 -56 -68087
rect 56 -67111 102 -67099
rect 56 -68087 62 -67111
rect 96 -68087 102 -67111
rect 56 -68099 102 -68087
rect -46 -68137 46 -68131
rect -46 -68171 -34 -68137
rect 34 -68171 46 -68137
rect -46 -68177 46 -68171
rect -46 -68245 46 -68239
rect -46 -68279 -34 -68245
rect 34 -68279 46 -68245
rect -46 -68285 46 -68279
rect -102 -68329 -56 -68317
rect -102 -69305 -96 -68329
rect -62 -69305 -56 -68329
rect -102 -69317 -56 -69305
rect 56 -68329 102 -68317
rect 56 -69305 62 -68329
rect 96 -69305 102 -68329
rect 56 -69317 102 -69305
rect -46 -69355 46 -69349
rect -46 -69389 -34 -69355
rect 34 -69389 46 -69355
rect -46 -69395 46 -69389
rect -46 -69463 46 -69457
rect -46 -69497 -34 -69463
rect 34 -69497 46 -69463
rect -46 -69503 46 -69497
rect -102 -69547 -56 -69535
rect -102 -70523 -96 -69547
rect -62 -70523 -56 -69547
rect -102 -70535 -56 -70523
rect 56 -69547 102 -69535
rect 56 -70523 62 -69547
rect 96 -70523 102 -69547
rect 56 -70535 102 -70523
rect -46 -70573 46 -70567
rect -46 -70607 -34 -70573
rect 34 -70607 46 -70573
rect -46 -70613 46 -70607
rect -46 -70681 46 -70675
rect -46 -70715 -34 -70681
rect 34 -70715 46 -70681
rect -46 -70721 46 -70715
rect -102 -70765 -56 -70753
rect -102 -71741 -96 -70765
rect -62 -71741 -56 -70765
rect -102 -71753 -56 -71741
rect 56 -70765 102 -70753
rect 56 -71741 62 -70765
rect 96 -71741 102 -70765
rect 56 -71753 102 -71741
rect -46 -71791 46 -71785
rect -46 -71825 -34 -71791
rect 34 -71825 46 -71791
rect -46 -71831 46 -71825
rect -46 -71899 46 -71893
rect -46 -71933 -34 -71899
rect 34 -71933 46 -71899
rect -46 -71939 46 -71933
rect -102 -71983 -56 -71971
rect -102 -72959 -96 -71983
rect -62 -72959 -56 -71983
rect -102 -72971 -56 -72959
rect 56 -71983 102 -71971
rect 56 -72959 62 -71983
rect 96 -72959 102 -71983
rect 56 -72971 102 -72959
rect -46 -73009 46 -73003
rect -46 -73043 -34 -73009
rect 34 -73043 46 -73009
rect -46 -73049 46 -73043
rect -46 -73117 46 -73111
rect -46 -73151 -34 -73117
rect 34 -73151 46 -73117
rect -46 -73157 46 -73151
rect -102 -73201 -56 -73189
rect -102 -74177 -96 -73201
rect -62 -74177 -56 -73201
rect -102 -74189 -56 -74177
rect 56 -73201 102 -73189
rect 56 -74177 62 -73201
rect 96 -74177 102 -73201
rect 56 -74189 102 -74177
rect -46 -74227 46 -74221
rect -46 -74261 -34 -74227
rect 34 -74261 46 -74227
rect -46 -74267 46 -74261
rect -46 -74335 46 -74329
rect -46 -74369 -34 -74335
rect 34 -74369 46 -74335
rect -46 -74375 46 -74369
rect -102 -74419 -56 -74407
rect -102 -75395 -96 -74419
rect -62 -75395 -56 -74419
rect -102 -75407 -56 -75395
rect 56 -74419 102 -74407
rect 56 -75395 62 -74419
rect 96 -75395 102 -74419
rect 56 -75407 102 -75395
rect -46 -75445 46 -75439
rect -46 -75479 -34 -75445
rect 34 -75479 46 -75445
rect -46 -75485 46 -75479
rect -46 -75553 46 -75547
rect -46 -75587 -34 -75553
rect 34 -75587 46 -75553
rect -46 -75593 46 -75587
rect -102 -75637 -56 -75625
rect -102 -76613 -96 -75637
rect -62 -76613 -56 -75637
rect -102 -76625 -56 -76613
rect 56 -75637 102 -75625
rect 56 -76613 62 -75637
rect 96 -76613 102 -75637
rect 56 -76625 102 -76613
rect -46 -76663 46 -76657
rect -46 -76697 -34 -76663
rect 34 -76697 46 -76663
rect -46 -76703 46 -76697
rect -46 -76771 46 -76765
rect -46 -76805 -34 -76771
rect 34 -76805 46 -76771
rect -46 -76811 46 -76805
rect -102 -76855 -56 -76843
rect -102 -77831 -96 -76855
rect -62 -77831 -56 -76855
rect -102 -77843 -56 -77831
rect 56 -76855 102 -76843
rect 56 -77831 62 -76855
rect 96 -77831 102 -76855
rect 56 -77843 102 -77831
rect -46 -77881 46 -77875
rect -46 -77915 -34 -77881
rect 34 -77915 46 -77881
rect -46 -77921 46 -77915
rect -46 -77989 46 -77983
rect -46 -78023 -34 -77989
rect 34 -78023 46 -77989
rect -46 -78029 46 -78023
rect -102 -78073 -56 -78061
rect -102 -79049 -96 -78073
rect -62 -79049 -56 -78073
rect -102 -79061 -56 -79049
rect 56 -78073 102 -78061
rect 56 -79049 62 -78073
rect 96 -79049 102 -78073
rect 56 -79061 102 -79049
rect -46 -79099 46 -79093
rect -46 -79133 -34 -79099
rect 34 -79133 46 -79099
rect -46 -79139 46 -79133
rect -46 -79207 46 -79201
rect -46 -79241 -34 -79207
rect 34 -79241 46 -79207
rect -46 -79247 46 -79241
rect -102 -79291 -56 -79279
rect -102 -80267 -96 -79291
rect -62 -80267 -56 -79291
rect -102 -80279 -56 -80267
rect 56 -79291 102 -79279
rect 56 -80267 62 -79291
rect 96 -80267 102 -79291
rect 56 -80279 102 -80267
rect -46 -80317 46 -80311
rect -46 -80351 -34 -80317
rect 34 -80351 46 -80317
rect -46 -80357 46 -80351
rect -46 -80425 46 -80419
rect -46 -80459 -34 -80425
rect 34 -80459 46 -80425
rect -46 -80465 46 -80459
rect -102 -80509 -56 -80497
rect -102 -81485 -96 -80509
rect -62 -81485 -56 -80509
rect -102 -81497 -56 -81485
rect 56 -80509 102 -80497
rect 56 -81485 62 -80509
rect 96 -81485 102 -80509
rect 56 -81497 102 -81485
rect -46 -81535 46 -81529
rect -46 -81569 -34 -81535
rect 34 -81569 46 -81535
rect -46 -81575 46 -81569
rect -46 -81643 46 -81637
rect -46 -81677 -34 -81643
rect 34 -81677 46 -81643
rect -46 -81683 46 -81677
rect -102 -81727 -56 -81715
rect -102 -82703 -96 -81727
rect -62 -82703 -56 -81727
rect -102 -82715 -56 -82703
rect 56 -81727 102 -81715
rect 56 -82703 62 -81727
rect 96 -82703 102 -81727
rect 56 -82715 102 -82703
rect -46 -82753 46 -82747
rect -46 -82787 -34 -82753
rect 34 -82787 46 -82753
rect -46 -82793 46 -82787
rect -46 -82861 46 -82855
rect -46 -82895 -34 -82861
rect 34 -82895 46 -82861
rect -46 -82901 46 -82895
rect -102 -82945 -56 -82933
rect -102 -83921 -96 -82945
rect -62 -83921 -56 -82945
rect -102 -83933 -56 -83921
rect 56 -82945 102 -82933
rect 56 -83921 62 -82945
rect 96 -83921 102 -82945
rect 56 -83933 102 -83921
rect -46 -83971 46 -83965
rect -46 -84005 -34 -83971
rect 34 -84005 46 -83971
rect -46 -84011 46 -84005
rect -46 -84079 46 -84073
rect -46 -84113 -34 -84079
rect 34 -84113 46 -84079
rect -46 -84119 46 -84113
rect -102 -84163 -56 -84151
rect -102 -85139 -96 -84163
rect -62 -85139 -56 -84163
rect -102 -85151 -56 -85139
rect 56 -84163 102 -84151
rect 56 -85139 62 -84163
rect 96 -85139 102 -84163
rect 56 -85151 102 -85139
rect -46 -85189 46 -85183
rect -46 -85223 -34 -85189
rect 34 -85223 46 -85189
rect -46 -85229 46 -85223
rect -46 -85297 46 -85291
rect -46 -85331 -34 -85297
rect 34 -85331 46 -85297
rect -46 -85337 46 -85331
rect -102 -85381 -56 -85369
rect -102 -86357 -96 -85381
rect -62 -86357 -56 -85381
rect -102 -86369 -56 -86357
rect 56 -85381 102 -85369
rect 56 -86357 62 -85381
rect 96 -86357 102 -85381
rect 56 -86369 102 -86357
rect -46 -86407 46 -86401
rect -46 -86441 -34 -86407
rect 34 -86441 46 -86407
rect -46 -86447 46 -86441
rect -46 -86515 46 -86509
rect -46 -86549 -34 -86515
rect 34 -86549 46 -86515
rect -46 -86555 46 -86549
rect -102 -86599 -56 -86587
rect -102 -87575 -96 -86599
rect -62 -87575 -56 -86599
rect -102 -87587 -56 -87575
rect 56 -86599 102 -86587
rect 56 -87575 62 -86599
rect 96 -87575 102 -86599
rect 56 -87587 102 -87575
rect -46 -87625 46 -87619
rect -46 -87659 -34 -87625
rect 34 -87659 46 -87625
rect -46 -87665 46 -87659
rect -46 -87733 46 -87727
rect -46 -87767 -34 -87733
rect 34 -87767 46 -87733
rect -46 -87773 46 -87767
rect -102 -87817 -56 -87805
rect -102 -88793 -96 -87817
rect -62 -88793 -56 -87817
rect -102 -88805 -56 -88793
rect 56 -87817 102 -87805
rect 56 -88793 62 -87817
rect 96 -88793 102 -87817
rect 56 -88805 102 -88793
rect -46 -88843 46 -88837
rect -46 -88877 -34 -88843
rect 34 -88877 46 -88843
rect -46 -88883 46 -88877
rect -46 -88951 46 -88945
rect -46 -88985 -34 -88951
rect 34 -88985 46 -88951
rect -46 -88991 46 -88985
rect -102 -89035 -56 -89023
rect -102 -90011 -96 -89035
rect -62 -90011 -56 -89035
rect -102 -90023 -56 -90011
rect 56 -89035 102 -89023
rect 56 -90011 62 -89035
rect 96 -90011 102 -89035
rect 56 -90023 102 -90011
rect -46 -90061 46 -90055
rect -46 -90095 -34 -90061
rect 34 -90095 46 -90061
rect -46 -90101 46 -90095
rect -46 -90169 46 -90163
rect -46 -90203 -34 -90169
rect 34 -90203 46 -90169
rect -46 -90209 46 -90203
rect -102 -90253 -56 -90241
rect -102 -91229 -96 -90253
rect -62 -91229 -56 -90253
rect -102 -91241 -56 -91229
rect 56 -90253 102 -90241
rect 56 -91229 62 -90253
rect 96 -91229 102 -90253
rect 56 -91241 102 -91229
rect -46 -91279 46 -91273
rect -46 -91313 -34 -91279
rect 34 -91313 46 -91279
rect -46 -91319 46 -91313
rect -46 -91387 46 -91381
rect -46 -91421 -34 -91387
rect 34 -91421 46 -91387
rect -46 -91427 46 -91421
rect -102 -91471 -56 -91459
rect -102 -92447 -96 -91471
rect -62 -92447 -56 -91471
rect -102 -92459 -56 -92447
rect 56 -91471 102 -91459
rect 56 -92447 62 -91471
rect 96 -92447 102 -91471
rect 56 -92459 102 -92447
rect -46 -92497 46 -92491
rect -46 -92531 -34 -92497
rect 34 -92531 46 -92497
rect -46 -92537 46 -92531
rect -46 -92605 46 -92599
rect -46 -92639 -34 -92605
rect 34 -92639 46 -92605
rect -46 -92645 46 -92639
rect -102 -92689 -56 -92677
rect -102 -93665 -96 -92689
rect -62 -93665 -56 -92689
rect -102 -93677 -56 -93665
rect 56 -92689 102 -92677
rect 56 -93665 62 -92689
rect 96 -93665 102 -92689
rect 56 -93677 102 -93665
rect -46 -93715 46 -93709
rect -46 -93749 -34 -93715
rect 34 -93749 46 -93715
rect -46 -93755 46 -93749
rect -46 -93823 46 -93817
rect -46 -93857 -34 -93823
rect 34 -93857 46 -93823
rect -46 -93863 46 -93857
rect -102 -93907 -56 -93895
rect -102 -94883 -96 -93907
rect -62 -94883 -56 -93907
rect -102 -94895 -56 -94883
rect 56 -93907 102 -93895
rect 56 -94883 62 -93907
rect 96 -94883 102 -93907
rect 56 -94895 102 -94883
rect -46 -94933 46 -94927
rect -46 -94967 -34 -94933
rect 34 -94967 46 -94933
rect -46 -94973 46 -94967
rect -46 -95041 46 -95035
rect -46 -95075 -34 -95041
rect 34 -95075 46 -95041
rect -46 -95081 46 -95075
rect -102 -95125 -56 -95113
rect -102 -96101 -96 -95125
rect -62 -96101 -56 -95125
rect -102 -96113 -56 -96101
rect 56 -95125 102 -95113
rect 56 -96101 62 -95125
rect 96 -96101 102 -95125
rect 56 -96113 102 -96101
rect -46 -96151 46 -96145
rect -46 -96185 -34 -96151
rect 34 -96185 46 -96151
rect -46 -96191 46 -96185
rect -46 -96259 46 -96253
rect -46 -96293 -34 -96259
rect 34 -96293 46 -96259
rect -46 -96299 46 -96293
rect -102 -96343 -56 -96331
rect -102 -97319 -96 -96343
rect -62 -97319 -56 -96343
rect -102 -97331 -56 -97319
rect 56 -96343 102 -96331
rect 56 -97319 62 -96343
rect 96 -97319 102 -96343
rect 56 -97331 102 -97319
rect -46 -97369 46 -97363
rect -46 -97403 -34 -97369
rect 34 -97403 46 -97369
rect -46 -97409 46 -97403
rect -46 -97477 46 -97471
rect -46 -97511 -34 -97477
rect 34 -97511 46 -97477
rect -46 -97517 46 -97511
rect -102 -97561 -56 -97549
rect -102 -98537 -96 -97561
rect -62 -98537 -56 -97561
rect -102 -98549 -56 -98537
rect 56 -97561 102 -97549
rect 56 -98537 62 -97561
rect 96 -98537 102 -97561
rect 56 -98549 102 -98537
rect -46 -98587 46 -98581
rect -46 -98621 -34 -98587
rect 34 -98621 46 -98587
rect -46 -98627 46 -98621
rect -46 -98695 46 -98689
rect -46 -98729 -34 -98695
rect 34 -98729 46 -98695
rect -46 -98735 46 -98729
rect -102 -98779 -56 -98767
rect -102 -99755 -96 -98779
rect -62 -99755 -56 -98779
rect -102 -99767 -56 -99755
rect 56 -98779 102 -98767
rect 56 -99755 62 -98779
rect 96 -99755 102 -98779
rect 56 -99767 102 -99755
rect -46 -99805 46 -99799
rect -46 -99839 -34 -99805
rect 34 -99839 46 -99805
rect -46 -99845 46 -99839
rect -46 -99913 46 -99907
rect -46 -99947 -34 -99913
rect 34 -99947 46 -99913
rect -46 -99953 46 -99947
rect -102 -99997 -56 -99985
rect -102 -100973 -96 -99997
rect -62 -100973 -56 -99997
rect -102 -100985 -56 -100973
rect 56 -99997 102 -99985
rect 56 -100973 62 -99997
rect 96 -100973 102 -99997
rect 56 -100985 102 -100973
rect -46 -101023 46 -101017
rect -46 -101057 -34 -101023
rect 34 -101057 46 -101023
rect -46 -101063 46 -101057
rect -46 -101131 46 -101125
rect -46 -101165 -34 -101131
rect 34 -101165 46 -101131
rect -46 -101171 46 -101165
rect -102 -101215 -56 -101203
rect -102 -102191 -96 -101215
rect -62 -102191 -56 -101215
rect -102 -102203 -56 -102191
rect 56 -101215 102 -101203
rect 56 -102191 62 -101215
rect 96 -102191 102 -101215
rect 56 -102203 102 -102191
rect -46 -102241 46 -102235
rect -46 -102275 -34 -102241
rect 34 -102275 46 -102241
rect -46 -102281 46 -102275
rect -46 -102349 46 -102343
rect -46 -102383 -34 -102349
rect 34 -102383 46 -102349
rect -46 -102389 46 -102383
rect -102 -102433 -56 -102421
rect -102 -103409 -96 -102433
rect -62 -103409 -56 -102433
rect -102 -103421 -56 -103409
rect 56 -102433 102 -102421
rect 56 -103409 62 -102433
rect 96 -103409 102 -102433
rect 56 -103421 102 -103409
rect -46 -103459 46 -103453
rect -46 -103493 -34 -103459
rect 34 -103493 46 -103459
rect -46 -103499 46 -103493
rect -46 -103567 46 -103561
rect -46 -103601 -34 -103567
rect 34 -103601 46 -103567
rect -46 -103607 46 -103601
rect -102 -103651 -56 -103639
rect -102 -104627 -96 -103651
rect -62 -104627 -56 -103651
rect -102 -104639 -56 -104627
rect 56 -103651 102 -103639
rect 56 -104627 62 -103651
rect 96 -104627 102 -103651
rect 56 -104639 102 -104627
rect -46 -104677 46 -104671
rect -46 -104711 -34 -104677
rect 34 -104711 46 -104677
rect -46 -104717 46 -104711
rect -46 -104785 46 -104779
rect -46 -104819 -34 -104785
rect 34 -104819 46 -104785
rect -46 -104825 46 -104819
rect -102 -104869 -56 -104857
rect -102 -105845 -96 -104869
rect -62 -105845 -56 -104869
rect -102 -105857 -56 -105845
rect 56 -104869 102 -104857
rect 56 -105845 62 -104869
rect 96 -105845 102 -104869
rect 56 -105857 102 -105845
rect -46 -105895 46 -105889
rect -46 -105929 -34 -105895
rect 34 -105929 46 -105895
rect -46 -105935 46 -105929
rect -46 -106003 46 -105997
rect -46 -106037 -34 -106003
rect 34 -106037 46 -106003
rect -46 -106043 46 -106037
rect -102 -106087 -56 -106075
rect -102 -107063 -96 -106087
rect -62 -107063 -56 -106087
rect -102 -107075 -56 -107063
rect 56 -106087 102 -106075
rect 56 -107063 62 -106087
rect 96 -107063 102 -106087
rect 56 -107075 102 -107063
rect -46 -107113 46 -107107
rect -46 -107147 -34 -107113
rect 34 -107147 46 -107113
rect -46 -107153 46 -107147
rect -46 -107221 46 -107215
rect -46 -107255 -34 -107221
rect 34 -107255 46 -107221
rect -46 -107261 46 -107255
rect -102 -107305 -56 -107293
rect -102 -108281 -96 -107305
rect -62 -108281 -56 -107305
rect -102 -108293 -56 -108281
rect 56 -107305 102 -107293
rect 56 -108281 62 -107305
rect 96 -108281 102 -107305
rect 56 -108293 102 -108281
rect -46 -108331 46 -108325
rect -46 -108365 -34 -108331
rect 34 -108365 46 -108331
rect -46 -108371 46 -108365
rect -46 -108439 46 -108433
rect -46 -108473 -34 -108439
rect 34 -108473 46 -108439
rect -46 -108479 46 -108473
rect -102 -108523 -56 -108511
rect -102 -109499 -96 -108523
rect -62 -109499 -56 -108523
rect -102 -109511 -56 -109499
rect 56 -108523 102 -108511
rect 56 -109499 62 -108523
rect 96 -109499 102 -108523
rect 56 -109511 102 -109499
rect -46 -109549 46 -109543
rect -46 -109583 -34 -109549
rect 34 -109583 46 -109549
rect -46 -109589 46 -109583
rect -46 -109657 46 -109651
rect -46 -109691 -34 -109657
rect 34 -109691 46 -109657
rect -46 -109697 46 -109691
rect -102 -109741 -56 -109729
rect -102 -110717 -96 -109741
rect -62 -110717 -56 -109741
rect -102 -110729 -56 -110717
rect 56 -109741 102 -109729
rect 56 -110717 62 -109741
rect 96 -110717 102 -109741
rect 56 -110729 102 -110717
rect -46 -110767 46 -110761
rect -46 -110801 -34 -110767
rect 34 -110801 46 -110767
rect -46 -110807 46 -110801
rect -46 -110875 46 -110869
rect -46 -110909 -34 -110875
rect 34 -110909 46 -110875
rect -46 -110915 46 -110909
rect -102 -110959 -56 -110947
rect -102 -111935 -96 -110959
rect -62 -111935 -56 -110959
rect -102 -111947 -56 -111935
rect 56 -110959 102 -110947
rect 56 -111935 62 -110959
rect 96 -111935 102 -110959
rect 56 -111947 102 -111935
rect -46 -111985 46 -111979
rect -46 -112019 -34 -111985
rect 34 -112019 46 -111985
rect -46 -112025 46 -112019
rect -46 -112093 46 -112087
rect -46 -112127 -34 -112093
rect 34 -112127 46 -112093
rect -46 -112133 46 -112127
rect -102 -112177 -56 -112165
rect -102 -113153 -96 -112177
rect -62 -113153 -56 -112177
rect -102 -113165 -56 -113153
rect 56 -112177 102 -112165
rect 56 -113153 62 -112177
rect 96 -113153 102 -112177
rect 56 -113165 102 -113153
rect -46 -113203 46 -113197
rect -46 -113237 -34 -113203
rect 34 -113237 46 -113203
rect -46 -113243 46 -113237
rect -46 -113311 46 -113305
rect -46 -113345 -34 -113311
rect 34 -113345 46 -113311
rect -46 -113351 46 -113345
rect -102 -113395 -56 -113383
rect -102 -114371 -96 -113395
rect -62 -114371 -56 -113395
rect -102 -114383 -56 -114371
rect 56 -113395 102 -113383
rect 56 -114371 62 -113395
rect 96 -114371 102 -113395
rect 56 -114383 102 -114371
rect -46 -114421 46 -114415
rect -46 -114455 -34 -114421
rect 34 -114455 46 -114421
rect -46 -114461 46 -114455
rect -46 -114529 46 -114523
rect -46 -114563 -34 -114529
rect 34 -114563 46 -114529
rect -46 -114569 46 -114563
rect -102 -114613 -56 -114601
rect -102 -115589 -96 -114613
rect -62 -115589 -56 -114613
rect -102 -115601 -56 -115589
rect 56 -114613 102 -114601
rect 56 -115589 62 -114613
rect 96 -115589 102 -114613
rect 56 -115601 102 -115589
rect -46 -115639 46 -115633
rect -46 -115673 -34 -115639
rect 34 -115673 46 -115639
rect -46 -115679 46 -115673
rect -46 -115747 46 -115741
rect -46 -115781 -34 -115747
rect 34 -115781 46 -115747
rect -46 -115787 46 -115781
rect -102 -115831 -56 -115819
rect -102 -116807 -96 -115831
rect -62 -116807 -56 -115831
rect -102 -116819 -56 -116807
rect 56 -115831 102 -115819
rect 56 -116807 62 -115831
rect 96 -116807 102 -115831
rect 56 -116819 102 -116807
rect -46 -116857 46 -116851
rect -46 -116891 -34 -116857
rect 34 -116891 46 -116857
rect -46 -116897 46 -116891
rect -46 -116965 46 -116959
rect -46 -116999 -34 -116965
rect 34 -116999 46 -116965
rect -46 -117005 46 -116999
rect -102 -117049 -56 -117037
rect -102 -118025 -96 -117049
rect -62 -118025 -56 -117049
rect -102 -118037 -56 -118025
rect 56 -117049 102 -117037
rect 56 -118025 62 -117049
rect 96 -118025 102 -117049
rect 56 -118037 102 -118025
rect -46 -118075 46 -118069
rect -46 -118109 -34 -118075
rect 34 -118109 46 -118075
rect -46 -118115 46 -118109
rect -46 -118183 46 -118177
rect -46 -118217 -34 -118183
rect 34 -118217 46 -118183
rect -46 -118223 46 -118217
rect -102 -118267 -56 -118255
rect -102 -119243 -96 -118267
rect -62 -119243 -56 -118267
rect -102 -119255 -56 -119243
rect 56 -118267 102 -118255
rect 56 -119243 62 -118267
rect 96 -119243 102 -118267
rect 56 -119255 102 -119243
rect -46 -119293 46 -119287
rect -46 -119327 -34 -119293
rect 34 -119327 46 -119293
rect -46 -119333 46 -119327
rect -46 -119401 46 -119395
rect -46 -119435 -34 -119401
rect 34 -119435 46 -119401
rect -46 -119441 46 -119435
rect -102 -119485 -56 -119473
rect -102 -120461 -96 -119485
rect -62 -120461 -56 -119485
rect -102 -120473 -56 -120461
rect 56 -119485 102 -119473
rect 56 -120461 62 -119485
rect 96 -120461 102 -119485
rect 56 -120473 102 -120461
rect -46 -120511 46 -120505
rect -46 -120545 -34 -120511
rect 34 -120545 46 -120511
rect -46 -120551 46 -120545
rect -46 -120619 46 -120613
rect -46 -120653 -34 -120619
rect 34 -120653 46 -120619
rect -46 -120659 46 -120653
rect -102 -120703 -56 -120691
rect -102 -121679 -96 -120703
rect -62 -121679 -56 -120703
rect -102 -121691 -56 -121679
rect 56 -120703 102 -120691
rect 56 -121679 62 -120703
rect 96 -121679 102 -120703
rect 56 -121691 102 -121679
rect -46 -121729 46 -121723
rect -46 -121763 -34 -121729
rect 34 -121763 46 -121729
rect -46 -121769 46 -121763
rect -46 -121837 46 -121831
rect -46 -121871 -34 -121837
rect 34 -121871 46 -121837
rect -46 -121877 46 -121871
rect -102 -121921 -56 -121909
rect -102 -122897 -96 -121921
rect -62 -122897 -56 -121921
rect -102 -122909 -56 -122897
rect 56 -121921 102 -121909
rect 56 -122897 62 -121921
rect 96 -122897 102 -121921
rect 56 -122909 102 -122897
rect -46 -122947 46 -122941
rect -46 -122981 -34 -122947
rect 34 -122981 46 -122947
rect -46 -122987 46 -122981
rect -46 -123055 46 -123049
rect -46 -123089 -34 -123055
rect 34 -123089 46 -123055
rect -46 -123095 46 -123089
rect -102 -123139 -56 -123127
rect -102 -124115 -96 -123139
rect -62 -124115 -56 -123139
rect -102 -124127 -56 -124115
rect 56 -123139 102 -123127
rect 56 -124115 62 -123139
rect 96 -124115 102 -123139
rect 56 -124127 102 -124115
rect -46 -124165 46 -124159
rect -46 -124199 -34 -124165
rect 34 -124199 46 -124165
rect -46 -124205 46 -124199
rect -46 -124273 46 -124267
rect -46 -124307 -34 -124273
rect 34 -124307 46 -124273
rect -46 -124313 46 -124307
rect -102 -124357 -56 -124345
rect -102 -125333 -96 -124357
rect -62 -125333 -56 -124357
rect -102 -125345 -56 -125333
rect 56 -124357 102 -124345
rect 56 -125333 62 -124357
rect 96 -125333 102 -124357
rect 56 -125345 102 -125333
rect -46 -125383 46 -125377
rect -46 -125417 -34 -125383
rect 34 -125417 46 -125383
rect -46 -125423 46 -125417
rect -46 -125491 46 -125485
rect -46 -125525 -34 -125491
rect 34 -125525 46 -125491
rect -46 -125531 46 -125525
rect -102 -125575 -56 -125563
rect -102 -126551 -96 -125575
rect -62 -126551 -56 -125575
rect -102 -126563 -56 -126551
rect 56 -125575 102 -125563
rect 56 -126551 62 -125575
rect 96 -126551 102 -125575
rect 56 -126563 102 -126551
rect -46 -126601 46 -126595
rect -46 -126635 -34 -126601
rect 34 -126635 46 -126601
rect -46 -126641 46 -126635
rect -46 -126709 46 -126703
rect -46 -126743 -34 -126709
rect 34 -126743 46 -126709
rect -46 -126749 46 -126743
rect -102 -126793 -56 -126781
rect -102 -127769 -96 -126793
rect -62 -127769 -56 -126793
rect -102 -127781 -56 -127769
rect 56 -126793 102 -126781
rect 56 -127769 62 -126793
rect 96 -127769 102 -126793
rect 56 -127781 102 -127769
rect -46 -127819 46 -127813
rect -46 -127853 -34 -127819
rect 34 -127853 46 -127819
rect -46 -127859 46 -127853
rect -46 -127927 46 -127921
rect -46 -127961 -34 -127927
rect 34 -127961 46 -127927
rect -46 -127967 46 -127961
rect -102 -128011 -56 -127999
rect -102 -128987 -96 -128011
rect -62 -128987 -56 -128011
rect -102 -128999 -56 -128987
rect 56 -128011 102 -127999
rect 56 -128987 62 -128011
rect 96 -128987 102 -128011
rect 56 -128999 102 -128987
rect -46 -129037 46 -129031
rect -46 -129071 -34 -129037
rect 34 -129071 46 -129037
rect -46 -129077 46 -129071
rect -46 -129145 46 -129139
rect -46 -129179 -34 -129145
rect 34 -129179 46 -129145
rect -46 -129185 46 -129179
rect -102 -129229 -56 -129217
rect -102 -130205 -96 -129229
rect -62 -130205 -56 -129229
rect -102 -130217 -56 -130205
rect 56 -129229 102 -129217
rect 56 -130205 62 -129229
rect 96 -130205 102 -129229
rect 56 -130217 102 -130205
rect -46 -130255 46 -130249
rect -46 -130289 -34 -130255
rect 34 -130289 46 -130255
rect -46 -130295 46 -130289
rect -46 -130363 46 -130357
rect -46 -130397 -34 -130363
rect 34 -130397 46 -130363
rect -46 -130403 46 -130397
rect -102 -130447 -56 -130435
rect -102 -131423 -96 -130447
rect -62 -131423 -56 -130447
rect -102 -131435 -56 -131423
rect 56 -130447 102 -130435
rect 56 -131423 62 -130447
rect 96 -131423 102 -130447
rect 56 -131435 102 -131423
rect -46 -131473 46 -131467
rect -46 -131507 -34 -131473
rect 34 -131507 46 -131473
rect -46 -131513 46 -131507
rect -46 -131581 46 -131575
rect -46 -131615 -34 -131581
rect 34 -131615 46 -131581
rect -46 -131621 46 -131615
rect -102 -131665 -56 -131653
rect -102 -132641 -96 -131665
rect -62 -132641 -56 -131665
rect -102 -132653 -56 -132641
rect 56 -131665 102 -131653
rect 56 -132641 62 -131665
rect 96 -132641 102 -131665
rect 56 -132653 102 -132641
rect -46 -132691 46 -132685
rect -46 -132725 -34 -132691
rect 34 -132725 46 -132691
rect -46 -132731 46 -132725
rect -46 -132799 46 -132793
rect -46 -132833 -34 -132799
rect 34 -132833 46 -132799
rect -46 -132839 46 -132833
rect -102 -132883 -56 -132871
rect -102 -133859 -96 -132883
rect -62 -133859 -56 -132883
rect -102 -133871 -56 -133859
rect 56 -132883 102 -132871
rect 56 -133859 62 -132883
rect 96 -133859 102 -132883
rect 56 -133871 102 -133859
rect -46 -133909 46 -133903
rect -46 -133943 -34 -133909
rect 34 -133943 46 -133909
rect -46 -133949 46 -133943
rect -46 -134017 46 -134011
rect -46 -134051 -34 -134017
rect 34 -134051 46 -134017
rect -46 -134057 46 -134051
rect -102 -134101 -56 -134089
rect -102 -135077 -96 -134101
rect -62 -135077 -56 -134101
rect -102 -135089 -56 -135077
rect 56 -134101 102 -134089
rect 56 -135077 62 -134101
rect 96 -135077 102 -134101
rect 56 -135089 102 -135077
rect -46 -135127 46 -135121
rect -46 -135161 -34 -135127
rect 34 -135161 46 -135127
rect -46 -135167 46 -135161
rect -46 -135235 46 -135229
rect -46 -135269 -34 -135235
rect 34 -135269 46 -135235
rect -46 -135275 46 -135269
rect -102 -135319 -56 -135307
rect -102 -136295 -96 -135319
rect -62 -136295 -56 -135319
rect -102 -136307 -56 -136295
rect 56 -135319 102 -135307
rect 56 -136295 62 -135319
rect 96 -136295 102 -135319
rect 56 -136307 102 -136295
rect -46 -136345 46 -136339
rect -46 -136379 -34 -136345
rect 34 -136379 46 -136345
rect -46 -136385 46 -136379
rect -46 -136453 46 -136447
rect -46 -136487 -34 -136453
rect 34 -136487 46 -136453
rect -46 -136493 46 -136487
rect -102 -136537 -56 -136525
rect -102 -137513 -96 -136537
rect -62 -137513 -56 -136537
rect -102 -137525 -56 -137513
rect 56 -136537 102 -136525
rect 56 -137513 62 -136537
rect 96 -137513 102 -136537
rect 56 -137525 102 -137513
rect -46 -137563 46 -137557
rect -46 -137597 -34 -137563
rect 34 -137597 46 -137563
rect -46 -137603 46 -137597
rect -46 -137671 46 -137665
rect -46 -137705 -34 -137671
rect 34 -137705 46 -137671
rect -46 -137711 46 -137705
rect -102 -137755 -56 -137743
rect -102 -138731 -96 -137755
rect -62 -138731 -56 -137755
rect -102 -138743 -56 -138731
rect 56 -137755 102 -137743
rect 56 -138731 62 -137755
rect 96 -138731 102 -137755
rect 56 -138743 102 -138731
rect -46 -138781 46 -138775
rect -46 -138815 -34 -138781
rect 34 -138815 46 -138781
rect -46 -138821 46 -138815
rect -46 -138889 46 -138883
rect -46 -138923 -34 -138889
rect 34 -138923 46 -138889
rect -46 -138929 46 -138923
rect -102 -138973 -56 -138961
rect -102 -139949 -96 -138973
rect -62 -139949 -56 -138973
rect -102 -139961 -56 -139949
rect 56 -138973 102 -138961
rect 56 -139949 62 -138973
rect 96 -139949 102 -138973
rect 56 -139961 102 -139949
rect -46 -139999 46 -139993
rect -46 -140033 -34 -139999
rect 34 -140033 46 -139999
rect -46 -140039 46 -140033
rect -46 -140107 46 -140101
rect -46 -140141 -34 -140107
rect 34 -140141 46 -140107
rect -46 -140147 46 -140141
rect -102 -140191 -56 -140179
rect -102 -141167 -96 -140191
rect -62 -141167 -56 -140191
rect -102 -141179 -56 -141167
rect 56 -140191 102 -140179
rect 56 -141167 62 -140191
rect 96 -141167 102 -140191
rect 56 -141179 102 -141167
rect -46 -141217 46 -141211
rect -46 -141251 -34 -141217
rect 34 -141251 46 -141217
rect -46 -141257 46 -141251
rect -46 -141325 46 -141319
rect -46 -141359 -34 -141325
rect 34 -141359 46 -141325
rect -46 -141365 46 -141359
rect -102 -141409 -56 -141397
rect -102 -142385 -96 -141409
rect -62 -142385 -56 -141409
rect -102 -142397 -56 -142385
rect 56 -141409 102 -141397
rect 56 -142385 62 -141409
rect 96 -142385 102 -141409
rect 56 -142397 102 -142385
rect -46 -142435 46 -142429
rect -46 -142469 -34 -142435
rect 34 -142469 46 -142435
rect -46 -142475 46 -142469
rect -46 -142543 46 -142537
rect -46 -142577 -34 -142543
rect 34 -142577 46 -142543
rect -46 -142583 46 -142577
rect -102 -142627 -56 -142615
rect -102 -143603 -96 -142627
rect -62 -143603 -56 -142627
rect -102 -143615 -56 -143603
rect 56 -142627 102 -142615
rect 56 -143603 62 -142627
rect 96 -143603 102 -142627
rect 56 -143615 102 -143603
rect -46 -143653 46 -143647
rect -46 -143687 -34 -143653
rect 34 -143687 46 -143653
rect -46 -143693 46 -143687
rect -46 -143761 46 -143755
rect -46 -143795 -34 -143761
rect 34 -143795 46 -143761
rect -46 -143801 46 -143795
rect -102 -143845 -56 -143833
rect -102 -144821 -96 -143845
rect -62 -144821 -56 -143845
rect -102 -144833 -56 -144821
rect 56 -143845 102 -143833
rect 56 -144821 62 -143845
rect 96 -144821 102 -143845
rect 56 -144833 102 -144821
rect -46 -144871 46 -144865
rect -46 -144905 -34 -144871
rect 34 -144905 46 -144871
rect -46 -144911 46 -144905
rect -46 -144979 46 -144973
rect -46 -145013 -34 -144979
rect 34 -145013 46 -144979
rect -46 -145019 46 -145013
rect -102 -145063 -56 -145051
rect -102 -146039 -96 -145063
rect -62 -146039 -56 -145063
rect -102 -146051 -56 -146039
rect 56 -145063 102 -145051
rect 56 -146039 62 -145063
rect 96 -146039 102 -145063
rect 56 -146051 102 -146039
rect -46 -146089 46 -146083
rect -46 -146123 -34 -146089
rect 34 -146123 46 -146089
rect -46 -146129 46 -146123
rect -46 -146197 46 -146191
rect -46 -146231 -34 -146197
rect 34 -146231 46 -146197
rect -46 -146237 46 -146231
rect -102 -146281 -56 -146269
rect -102 -147257 -96 -146281
rect -62 -147257 -56 -146281
rect -102 -147269 -56 -147257
rect 56 -146281 102 -146269
rect 56 -147257 62 -146281
rect 96 -147257 102 -146281
rect 56 -147269 102 -147257
rect -46 -147307 46 -147301
rect -46 -147341 -34 -147307
rect 34 -147341 46 -147307
rect -46 -147347 46 -147341
rect -46 -147415 46 -147409
rect -46 -147449 -34 -147415
rect 34 -147449 46 -147415
rect -46 -147455 46 -147449
rect -102 -147499 -56 -147487
rect -102 -148475 -96 -147499
rect -62 -148475 -56 -147499
rect -102 -148487 -56 -148475
rect 56 -147499 102 -147487
rect 56 -148475 62 -147499
rect 96 -148475 102 -147499
rect 56 -148487 102 -148475
rect -46 -148525 46 -148519
rect -46 -148559 -34 -148525
rect 34 -148559 46 -148525
rect -46 -148565 46 -148559
rect -46 -148633 46 -148627
rect -46 -148667 -34 -148633
rect 34 -148667 46 -148633
rect -46 -148673 46 -148667
rect -102 -148717 -56 -148705
rect -102 -149693 -96 -148717
rect -62 -149693 -56 -148717
rect -102 -149705 -56 -149693
rect 56 -148717 102 -148705
rect 56 -149693 62 -148717
rect 96 -149693 102 -148717
rect 56 -149705 102 -149693
rect -46 -149743 46 -149737
rect -46 -149777 -34 -149743
rect 34 -149777 46 -149743
rect -46 -149783 46 -149777
rect -46 -149851 46 -149845
rect -46 -149885 -34 -149851
rect 34 -149885 46 -149851
rect -46 -149891 46 -149885
rect -102 -149935 -56 -149923
rect -102 -150911 -96 -149935
rect -62 -150911 -56 -149935
rect -102 -150923 -56 -150911
rect 56 -149935 102 -149923
rect 56 -150911 62 -149935
rect 96 -150911 102 -149935
rect 56 -150923 102 -150911
rect -46 -150961 46 -150955
rect -46 -150995 -34 -150961
rect 34 -150995 46 -150961
rect -46 -151001 46 -150995
rect -46 -151069 46 -151063
rect -46 -151103 -34 -151069
rect 34 -151103 46 -151069
rect -46 -151109 46 -151103
rect -102 -151153 -56 -151141
rect -102 -152129 -96 -151153
rect -62 -152129 -56 -151153
rect -102 -152141 -56 -152129
rect 56 -151153 102 -151141
rect 56 -152129 62 -151153
rect 96 -152129 102 -151153
rect 56 -152141 102 -152129
rect -46 -152179 46 -152173
rect -46 -152213 -34 -152179
rect 34 -152213 46 -152179
rect -46 -152219 46 -152213
rect -46 -152287 46 -152281
rect -46 -152321 -34 -152287
rect 34 -152321 46 -152287
rect -46 -152327 46 -152321
rect -102 -152371 -56 -152359
rect -102 -153347 -96 -152371
rect -62 -153347 -56 -152371
rect -102 -153359 -56 -153347
rect 56 -152371 102 -152359
rect 56 -153347 62 -152371
rect 96 -153347 102 -152371
rect 56 -153359 102 -153347
rect -46 -153397 46 -153391
rect -46 -153431 -34 -153397
rect 34 -153431 46 -153397
rect -46 -153437 46 -153431
rect -46 -153505 46 -153499
rect -46 -153539 -34 -153505
rect 34 -153539 46 -153505
rect -46 -153545 46 -153539
rect -102 -153589 -56 -153577
rect -102 -154565 -96 -153589
rect -62 -154565 -56 -153589
rect -102 -154577 -56 -154565
rect 56 -153589 102 -153577
rect 56 -154565 62 -153589
rect 96 -154565 102 -153589
rect 56 -154577 102 -154565
rect -46 -154615 46 -154609
rect -46 -154649 -34 -154615
rect 34 -154649 46 -154615
rect -46 -154655 46 -154649
rect -46 -154723 46 -154717
rect -46 -154757 -34 -154723
rect 34 -154757 46 -154723
rect -46 -154763 46 -154757
rect -102 -154807 -56 -154795
rect -102 -155783 -96 -154807
rect -62 -155783 -56 -154807
rect -102 -155795 -56 -155783
rect 56 -154807 102 -154795
rect 56 -155783 62 -154807
rect 96 -155783 102 -154807
rect 56 -155795 102 -155783
rect -46 -155833 46 -155827
rect -46 -155867 -34 -155833
rect 34 -155867 46 -155833
rect -46 -155873 46 -155867
rect -46 -155941 46 -155935
rect -46 -155975 -34 -155941
rect 34 -155975 46 -155941
rect -46 -155981 46 -155975
rect -102 -156025 -56 -156013
rect -102 -157001 -96 -156025
rect -62 -157001 -56 -156025
rect -102 -157013 -56 -157001
rect 56 -156025 102 -156013
rect 56 -157001 62 -156025
rect 96 -157001 102 -156025
rect 56 -157013 102 -157001
rect -46 -157051 46 -157045
rect -46 -157085 -34 -157051
rect 34 -157085 46 -157051
rect -46 -157091 46 -157085
rect -46 -157159 46 -157153
rect -46 -157193 -34 -157159
rect 34 -157193 46 -157159
rect -46 -157199 46 -157193
rect -102 -157243 -56 -157231
rect -102 -158219 -96 -157243
rect -62 -158219 -56 -157243
rect -102 -158231 -56 -158219
rect 56 -157243 102 -157231
rect 56 -158219 62 -157243
rect 96 -158219 102 -157243
rect 56 -158231 102 -158219
rect -46 -158269 46 -158263
rect -46 -158303 -34 -158269
rect 34 -158303 46 -158269
rect -46 -158309 46 -158303
rect -46 -158377 46 -158371
rect -46 -158411 -34 -158377
rect 34 -158411 46 -158377
rect -46 -158417 46 -158411
rect -102 -158461 -56 -158449
rect -102 -159437 -96 -158461
rect -62 -159437 -56 -158461
rect -102 -159449 -56 -159437
rect 56 -158461 102 -158449
rect 56 -159437 62 -158461
rect 96 -159437 102 -158461
rect 56 -159449 102 -159437
rect -46 -159487 46 -159481
rect -46 -159521 -34 -159487
rect 34 -159521 46 -159487
rect -46 -159527 46 -159521
rect -46 -159595 46 -159589
rect -46 -159629 -34 -159595
rect 34 -159629 46 -159595
rect -46 -159635 46 -159629
rect -102 -159679 -56 -159667
rect -102 -160655 -96 -159679
rect -62 -160655 -56 -159679
rect -102 -160667 -56 -160655
rect 56 -159679 102 -159667
rect 56 -160655 62 -159679
rect 96 -160655 102 -159679
rect 56 -160667 102 -160655
rect -46 -160705 46 -160699
rect -46 -160739 -34 -160705
rect 34 -160739 46 -160705
rect -46 -160745 46 -160739
rect -46 -160813 46 -160807
rect -46 -160847 -34 -160813
rect 34 -160847 46 -160813
rect -46 -160853 46 -160847
rect -102 -160897 -56 -160885
rect -102 -161873 -96 -160897
rect -62 -161873 -56 -160897
rect -102 -161885 -56 -161873
rect 56 -160897 102 -160885
rect 56 -161873 62 -160897
rect 96 -161873 102 -160897
rect 56 -161885 102 -161873
rect -46 -161923 46 -161917
rect -46 -161957 -34 -161923
rect 34 -161957 46 -161923
rect -46 -161963 46 -161957
rect -46 -162031 46 -162025
rect -46 -162065 -34 -162031
rect 34 -162065 46 -162031
rect -46 -162071 46 -162065
rect -102 -162115 -56 -162103
rect -102 -163091 -96 -162115
rect -62 -163091 -56 -162115
rect -102 -163103 -56 -163091
rect 56 -162115 102 -162103
rect 56 -163091 62 -162115
rect 96 -163091 102 -162115
rect 56 -163103 102 -163091
rect -46 -163141 46 -163135
rect -46 -163175 -34 -163141
rect 34 -163175 46 -163141
rect -46 -163181 46 -163175
rect -46 -163249 46 -163243
rect -46 -163283 -34 -163249
rect 34 -163283 46 -163249
rect -46 -163289 46 -163283
rect -102 -163333 -56 -163321
rect -102 -164309 -96 -163333
rect -62 -164309 -56 -163333
rect -102 -164321 -56 -164309
rect 56 -163333 102 -163321
rect 56 -164309 62 -163333
rect 96 -164309 102 -163333
rect 56 -164321 102 -164309
rect -46 -164359 46 -164353
rect -46 -164393 -34 -164359
rect 34 -164393 46 -164359
rect -46 -164399 46 -164393
rect -46 -164467 46 -164461
rect -46 -164501 -34 -164467
rect 34 -164501 46 -164467
rect -46 -164507 46 -164501
rect -102 -164551 -56 -164539
rect -102 -165527 -96 -164551
rect -62 -165527 -56 -164551
rect -102 -165539 -56 -165527
rect 56 -164551 102 -164539
rect 56 -165527 62 -164551
rect 96 -165527 102 -164551
rect 56 -165539 102 -165527
rect -46 -165577 46 -165571
rect -46 -165611 -34 -165577
rect 34 -165611 46 -165577
rect -46 -165617 46 -165611
rect -46 -165685 46 -165679
rect -46 -165719 -34 -165685
rect 34 -165719 46 -165685
rect -46 -165725 46 -165719
rect -102 -165769 -56 -165757
rect -102 -166745 -96 -165769
rect -62 -166745 -56 -165769
rect -102 -166757 -56 -166745
rect 56 -165769 102 -165757
rect 56 -166745 62 -165769
rect 96 -166745 102 -165769
rect 56 -166757 102 -166745
rect -46 -166795 46 -166789
rect -46 -166829 -34 -166795
rect 34 -166829 46 -166795
rect -46 -166835 46 -166829
rect -46 -166903 46 -166897
rect -46 -166937 -34 -166903
rect 34 -166937 46 -166903
rect -46 -166943 46 -166937
rect -102 -166987 -56 -166975
rect -102 -167963 -96 -166987
rect -62 -167963 -56 -166987
rect -102 -167975 -56 -167963
rect 56 -166987 102 -166975
rect 56 -167963 62 -166987
rect 96 -167963 102 -166987
rect 56 -167975 102 -167963
rect -46 -168013 46 -168007
rect -46 -168047 -34 -168013
rect 34 -168047 46 -168013
rect -46 -168053 46 -168047
rect -46 -168121 46 -168115
rect -46 -168155 -34 -168121
rect 34 -168155 46 -168121
rect -46 -168161 46 -168155
rect -102 -168205 -56 -168193
rect -102 -169181 -96 -168205
rect -62 -169181 -56 -168205
rect -102 -169193 -56 -169181
rect 56 -168205 102 -168193
rect 56 -169181 62 -168205
rect 96 -169181 102 -168205
rect 56 -169193 102 -169181
rect -46 -169231 46 -169225
rect -46 -169265 -34 -169231
rect 34 -169265 46 -169231
rect -46 -169271 46 -169265
rect -46 -169339 46 -169333
rect -46 -169373 -34 -169339
rect 34 -169373 46 -169339
rect -46 -169379 46 -169373
rect -102 -169423 -56 -169411
rect -102 -170399 -96 -169423
rect -62 -170399 -56 -169423
rect -102 -170411 -56 -170399
rect 56 -169423 102 -169411
rect 56 -170399 62 -169423
rect 96 -170399 102 -169423
rect 56 -170411 102 -170399
rect -46 -170449 46 -170443
rect -46 -170483 -34 -170449
rect 34 -170483 46 -170449
rect -46 -170489 46 -170483
rect -46 -170557 46 -170551
rect -46 -170591 -34 -170557
rect 34 -170591 46 -170557
rect -46 -170597 46 -170591
rect -102 -170641 -56 -170629
rect -102 -171617 -96 -170641
rect -62 -171617 -56 -170641
rect -102 -171629 -56 -171617
rect 56 -170641 102 -170629
rect 56 -171617 62 -170641
rect 96 -171617 102 -170641
rect 56 -171629 102 -171617
rect -46 -171667 46 -171661
rect -46 -171701 -34 -171667
rect 34 -171701 46 -171667
rect -46 -171707 46 -171701
rect -46 -171775 46 -171769
rect -46 -171809 -34 -171775
rect 34 -171809 46 -171775
rect -46 -171815 46 -171809
rect -102 -171859 -56 -171847
rect -102 -172835 -96 -171859
rect -62 -172835 -56 -171859
rect -102 -172847 -56 -172835
rect 56 -171859 102 -171847
rect 56 -172835 62 -171859
rect 96 -172835 102 -171859
rect 56 -172847 102 -172835
rect -46 -172885 46 -172879
rect -46 -172919 -34 -172885
rect 34 -172919 46 -172885
rect -46 -172925 46 -172919
rect -46 -172993 46 -172987
rect -46 -173027 -34 -172993
rect 34 -173027 46 -172993
rect -46 -173033 46 -173027
rect -102 -173077 -56 -173065
rect -102 -174053 -96 -173077
rect -62 -174053 -56 -173077
rect -102 -174065 -56 -174053
rect 56 -173077 102 -173065
rect 56 -174053 62 -173077
rect 96 -174053 102 -173077
rect 56 -174065 102 -174053
rect -46 -174103 46 -174097
rect -46 -174137 -34 -174103
rect 34 -174137 46 -174103
rect -46 -174143 46 -174137
rect -46 -174211 46 -174205
rect -46 -174245 -34 -174211
rect 34 -174245 46 -174211
rect -46 -174251 46 -174245
rect -102 -174295 -56 -174283
rect -102 -175271 -96 -174295
rect -62 -175271 -56 -174295
rect -102 -175283 -56 -175271
rect 56 -174295 102 -174283
rect 56 -175271 62 -174295
rect 96 -175271 102 -174295
rect 56 -175283 102 -175271
rect -46 -175321 46 -175315
rect -46 -175355 -34 -175321
rect 34 -175355 46 -175321
rect -46 -175361 46 -175355
rect -46 -175429 46 -175423
rect -46 -175463 -34 -175429
rect 34 -175463 46 -175429
rect -46 -175469 46 -175463
rect -102 -175513 -56 -175501
rect -102 -176489 -96 -175513
rect -62 -176489 -56 -175513
rect -102 -176501 -56 -176489
rect 56 -175513 102 -175501
rect 56 -176489 62 -175513
rect 96 -176489 102 -175513
rect 56 -176501 102 -176489
rect -46 -176539 46 -176533
rect -46 -176573 -34 -176539
rect 34 -176573 46 -176539
rect -46 -176579 46 -176573
rect -46 -176647 46 -176641
rect -46 -176681 -34 -176647
rect 34 -176681 46 -176647
rect -46 -176687 46 -176681
rect -102 -176731 -56 -176719
rect -102 -177707 -96 -176731
rect -62 -177707 -56 -176731
rect -102 -177719 -56 -177707
rect 56 -176731 102 -176719
rect 56 -177707 62 -176731
rect 96 -177707 102 -176731
rect 56 -177719 102 -177707
rect -46 -177757 46 -177751
rect -46 -177791 -34 -177757
rect 34 -177791 46 -177757
rect -46 -177797 46 -177791
rect -46 -177865 46 -177859
rect -46 -177899 -34 -177865
rect 34 -177899 46 -177865
rect -46 -177905 46 -177899
rect -102 -177949 -56 -177937
rect -102 -178925 -96 -177949
rect -62 -178925 -56 -177949
rect -102 -178937 -56 -178925
rect 56 -177949 102 -177937
rect 56 -178925 62 -177949
rect 96 -178925 102 -177949
rect 56 -178937 102 -178925
rect -46 -178975 46 -178969
rect -46 -179009 -34 -178975
rect 34 -179009 46 -178975
rect -46 -179015 46 -179009
rect -46 -179083 46 -179077
rect -46 -179117 -34 -179083
rect 34 -179117 46 -179083
rect -46 -179123 46 -179117
rect -102 -179167 -56 -179155
rect -102 -180143 -96 -179167
rect -62 -180143 -56 -179167
rect -102 -180155 -56 -180143
rect 56 -179167 102 -179155
rect 56 -180143 62 -179167
rect 96 -180143 102 -179167
rect 56 -180155 102 -180143
rect -46 -180193 46 -180187
rect -46 -180227 -34 -180193
rect 34 -180227 46 -180193
rect -46 -180233 46 -180227
rect -46 -180301 46 -180295
rect -46 -180335 -34 -180301
rect 34 -180335 46 -180301
rect -46 -180341 46 -180335
rect -102 -180385 -56 -180373
rect -102 -181361 -96 -180385
rect -62 -181361 -56 -180385
rect -102 -181373 -56 -181361
rect 56 -180385 102 -180373
rect 56 -181361 62 -180385
rect 96 -181361 102 -180385
rect 56 -181373 102 -181361
rect -46 -181411 46 -181405
rect -46 -181445 -34 -181411
rect 34 -181445 46 -181411
rect -46 -181451 46 -181445
rect -46 -181519 46 -181513
rect -46 -181553 -34 -181519
rect 34 -181553 46 -181519
rect -46 -181559 46 -181553
rect -102 -181603 -56 -181591
rect -102 -182579 -96 -181603
rect -62 -182579 -56 -181603
rect -102 -182591 -56 -182579
rect 56 -181603 102 -181591
rect 56 -182579 62 -181603
rect 96 -182579 102 -181603
rect 56 -182591 102 -182579
rect -46 -182629 46 -182623
rect -46 -182663 -34 -182629
rect 34 -182663 46 -182629
rect -46 -182669 46 -182663
rect -46 -182737 46 -182731
rect -46 -182771 -34 -182737
rect 34 -182771 46 -182737
rect -46 -182777 46 -182771
rect -102 -182821 -56 -182809
rect -102 -183797 -96 -182821
rect -62 -183797 -56 -182821
rect -102 -183809 -56 -183797
rect 56 -182821 102 -182809
rect 56 -183797 62 -182821
rect 96 -183797 102 -182821
rect 56 -183809 102 -183797
rect -46 -183847 46 -183841
rect -46 -183881 -34 -183847
rect 34 -183881 46 -183847
rect -46 -183887 46 -183881
rect -46 -183955 46 -183949
rect -46 -183989 -34 -183955
rect 34 -183989 46 -183955
rect -46 -183995 46 -183989
rect -102 -184039 -56 -184027
rect -102 -185015 -96 -184039
rect -62 -185015 -56 -184039
rect -102 -185027 -56 -185015
rect 56 -184039 102 -184027
rect 56 -185015 62 -184039
rect 96 -185015 102 -184039
rect 56 -185027 102 -185015
rect -46 -185065 46 -185059
rect -46 -185099 -34 -185065
rect 34 -185099 46 -185065
rect -46 -185105 46 -185099
rect -46 -185173 46 -185167
rect -46 -185207 -34 -185173
rect 34 -185207 46 -185173
rect -46 -185213 46 -185207
rect -102 -185257 -56 -185245
rect -102 -186233 -96 -185257
rect -62 -186233 -56 -185257
rect -102 -186245 -56 -186233
rect 56 -185257 102 -185245
rect 56 -186233 62 -185257
rect 96 -186233 102 -185257
rect 56 -186245 102 -186233
rect -46 -186283 46 -186277
rect -46 -186317 -34 -186283
rect 34 -186317 46 -186283
rect -46 -186323 46 -186317
rect -46 -186391 46 -186385
rect -46 -186425 -34 -186391
rect 34 -186425 46 -186391
rect -46 -186431 46 -186425
rect -102 -186475 -56 -186463
rect -102 -187451 -96 -186475
rect -62 -187451 -56 -186475
rect -102 -187463 -56 -187451
rect 56 -186475 102 -186463
rect 56 -187451 62 -186475
rect 96 -187451 102 -186475
rect 56 -187463 102 -187451
rect -46 -187501 46 -187495
rect -46 -187535 -34 -187501
rect 34 -187535 46 -187501
rect -46 -187541 46 -187535
rect -46 -187609 46 -187603
rect -46 -187643 -34 -187609
rect 34 -187643 46 -187609
rect -46 -187649 46 -187643
rect -102 -187693 -56 -187681
rect -102 -188669 -96 -187693
rect -62 -188669 -56 -187693
rect -102 -188681 -56 -188669
rect 56 -187693 102 -187681
rect 56 -188669 62 -187693
rect 96 -188669 102 -187693
rect 56 -188681 102 -188669
rect -46 -188719 46 -188713
rect -46 -188753 -34 -188719
rect 34 -188753 46 -188719
rect -46 -188759 46 -188753
rect -46 -188827 46 -188821
rect -46 -188861 -34 -188827
rect 34 -188861 46 -188827
rect -46 -188867 46 -188861
rect -102 -188911 -56 -188899
rect -102 -189887 -96 -188911
rect -62 -189887 -56 -188911
rect -102 -189899 -56 -189887
rect 56 -188911 102 -188899
rect 56 -189887 62 -188911
rect 96 -189887 102 -188911
rect 56 -189899 102 -189887
rect -46 -189937 46 -189931
rect -46 -189971 -34 -189937
rect 34 -189971 46 -189937
rect -46 -189977 46 -189971
rect -46 -190045 46 -190039
rect -46 -190079 -34 -190045
rect 34 -190079 46 -190045
rect -46 -190085 46 -190079
rect -102 -190129 -56 -190117
rect -102 -191105 -96 -190129
rect -62 -191105 -56 -190129
rect -102 -191117 -56 -191105
rect 56 -190129 102 -190117
rect 56 -191105 62 -190129
rect 96 -191105 102 -190129
rect 56 -191117 102 -191105
rect -46 -191155 46 -191149
rect -46 -191189 -34 -191155
rect 34 -191189 46 -191155
rect -46 -191195 46 -191189
rect -46 -191263 46 -191257
rect -46 -191297 -34 -191263
rect 34 -191297 46 -191263
rect -46 -191303 46 -191297
rect -102 -191347 -56 -191335
rect -102 -192323 -96 -191347
rect -62 -192323 -56 -191347
rect -102 -192335 -56 -192323
rect 56 -191347 102 -191335
rect 56 -192323 62 -191347
rect 96 -192323 102 -191347
rect 56 -192335 102 -192323
rect -46 -192373 46 -192367
rect -46 -192407 -34 -192373
rect 34 -192407 46 -192373
rect -46 -192413 46 -192407
rect -46 -192481 46 -192475
rect -46 -192515 -34 -192481
rect 34 -192515 46 -192481
rect -46 -192521 46 -192515
rect -102 -192565 -56 -192553
rect -102 -193541 -96 -192565
rect -62 -193541 -56 -192565
rect -102 -193553 -56 -193541
rect 56 -192565 102 -192553
rect 56 -193541 62 -192565
rect 96 -193541 102 -192565
rect 56 -193553 102 -193541
rect -46 -193591 46 -193585
rect -46 -193625 -34 -193591
rect 34 -193625 46 -193591
rect -46 -193631 46 -193625
rect -46 -193699 46 -193693
rect -46 -193733 -34 -193699
rect 34 -193733 46 -193699
rect -46 -193739 46 -193733
rect -102 -193783 -56 -193771
rect -102 -194759 -96 -193783
rect -62 -194759 -56 -193783
rect -102 -194771 -56 -194759
rect 56 -193783 102 -193771
rect 56 -194759 62 -193783
rect 96 -194759 102 -193783
rect 56 -194771 102 -194759
rect -46 -194809 46 -194803
rect -46 -194843 -34 -194809
rect 34 -194843 46 -194809
rect -46 -194849 46 -194843
rect -46 -194917 46 -194911
rect -46 -194951 -34 -194917
rect 34 -194951 46 -194917
rect -46 -194957 46 -194951
rect -102 -195001 -56 -194989
rect -102 -195977 -96 -195001
rect -62 -195977 -56 -195001
rect -102 -195989 -56 -195977
rect 56 -195001 102 -194989
rect 56 -195977 62 -195001
rect 96 -195977 102 -195001
rect 56 -195989 102 -195977
rect -46 -196027 46 -196021
rect -46 -196061 -34 -196027
rect 34 -196061 46 -196027
rect -46 -196067 46 -196061
rect -46 -196135 46 -196129
rect -46 -196169 -34 -196135
rect 34 -196169 46 -196135
rect -46 -196175 46 -196169
rect -102 -196219 -56 -196207
rect -102 -197195 -96 -196219
rect -62 -197195 -56 -196219
rect -102 -197207 -56 -197195
rect 56 -196219 102 -196207
rect 56 -197195 62 -196219
rect 96 -197195 102 -196219
rect 56 -197207 102 -197195
rect -46 -197245 46 -197239
rect -46 -197279 -34 -197245
rect 34 -197279 46 -197245
rect -46 -197285 46 -197279
rect -46 -197353 46 -197347
rect -46 -197387 -34 -197353
rect 34 -197387 46 -197353
rect -46 -197393 46 -197387
rect -102 -197437 -56 -197425
rect -102 -198413 -96 -197437
rect -62 -198413 -56 -197437
rect -102 -198425 -56 -198413
rect 56 -197437 102 -197425
rect 56 -198413 62 -197437
rect 96 -198413 102 -197437
rect 56 -198425 102 -198413
rect -46 -198463 46 -198457
rect -46 -198497 -34 -198463
rect 34 -198497 46 -198463
rect -46 -198503 46 -198497
rect -46 -198571 46 -198565
rect -46 -198605 -34 -198571
rect 34 -198605 46 -198571
rect -46 -198611 46 -198605
rect -102 -198655 -56 -198643
rect -102 -199631 -96 -198655
rect -62 -199631 -56 -198655
rect -102 -199643 -56 -199631
rect 56 -198655 102 -198643
rect 56 -199631 62 -198655
rect 96 -199631 102 -198655
rect 56 -199643 102 -199631
rect -46 -199681 46 -199675
rect -46 -199715 -34 -199681
rect 34 -199715 46 -199681
rect -46 -199721 46 -199715
rect -46 -199789 46 -199783
rect -46 -199823 -34 -199789
rect 34 -199823 46 -199789
rect -46 -199829 46 -199823
rect -102 -199873 -56 -199861
rect -102 -200849 -96 -199873
rect -62 -200849 -56 -199873
rect -102 -200861 -56 -200849
rect 56 -199873 102 -199861
rect 56 -200849 62 -199873
rect 96 -200849 102 -199873
rect 56 -200861 102 -200849
rect -46 -200899 46 -200893
rect -46 -200933 -34 -200899
rect 34 -200933 46 -200899
rect -46 -200939 46 -200933
rect -46 -201007 46 -201001
rect -46 -201041 -34 -201007
rect 34 -201041 46 -201007
rect -46 -201047 46 -201041
rect -102 -201091 -56 -201079
rect -102 -202067 -96 -201091
rect -62 -202067 -56 -201091
rect -102 -202079 -56 -202067
rect 56 -201091 102 -201079
rect 56 -202067 62 -201091
rect 96 -202067 102 -201091
rect 56 -202079 102 -202067
rect -46 -202117 46 -202111
rect -46 -202151 -34 -202117
rect 34 -202151 46 -202117
rect -46 -202157 46 -202151
rect -46 -202225 46 -202219
rect -46 -202259 -34 -202225
rect 34 -202259 46 -202225
rect -46 -202265 46 -202259
rect -102 -202309 -56 -202297
rect -102 -203285 -96 -202309
rect -62 -203285 -56 -202309
rect -102 -203297 -56 -203285
rect 56 -202309 102 -202297
rect 56 -203285 62 -202309
rect 96 -203285 102 -202309
rect 56 -203297 102 -203285
rect -46 -203335 46 -203329
rect -46 -203369 -34 -203335
rect 34 -203369 46 -203335
rect -46 -203375 46 -203369
rect -46 -203443 46 -203437
rect -46 -203477 -34 -203443
rect 34 -203477 46 -203443
rect -46 -203483 46 -203477
rect -102 -203527 -56 -203515
rect -102 -204503 -96 -203527
rect -62 -204503 -56 -203527
rect -102 -204515 -56 -204503
rect 56 -203527 102 -203515
rect 56 -204503 62 -203527
rect 96 -204503 102 -203527
rect 56 -204515 102 -204503
rect -46 -204553 46 -204547
rect -46 -204587 -34 -204553
rect 34 -204587 46 -204553
rect -46 -204593 46 -204587
rect -46 -204661 46 -204655
rect -46 -204695 -34 -204661
rect 34 -204695 46 -204661
rect -46 -204701 46 -204695
rect -102 -204745 -56 -204733
rect -102 -205721 -96 -204745
rect -62 -205721 -56 -204745
rect -102 -205733 -56 -205721
rect 56 -204745 102 -204733
rect 56 -205721 62 -204745
rect 96 -205721 102 -204745
rect 56 -205733 102 -205721
rect -46 -205771 46 -205765
rect -46 -205805 -34 -205771
rect 34 -205805 46 -205771
rect -46 -205811 46 -205805
rect -46 -205879 46 -205873
rect -46 -205913 -34 -205879
rect 34 -205913 46 -205879
rect -46 -205919 46 -205913
rect -102 -205963 -56 -205951
rect -102 -206939 -96 -205963
rect -62 -206939 -56 -205963
rect -102 -206951 -56 -206939
rect 56 -205963 102 -205951
rect 56 -206939 62 -205963
rect 96 -206939 102 -205963
rect 56 -206951 102 -206939
rect -46 -206989 46 -206983
rect -46 -207023 -34 -206989
rect 34 -207023 46 -206989
rect -46 -207029 46 -207023
rect -46 -207097 46 -207091
rect -46 -207131 -34 -207097
rect 34 -207131 46 -207097
rect -46 -207137 46 -207131
rect -102 -207181 -56 -207169
rect -102 -208157 -96 -207181
rect -62 -208157 -56 -207181
rect -102 -208169 -56 -208157
rect 56 -207181 102 -207169
rect 56 -208157 62 -207181
rect 96 -208157 102 -207181
rect 56 -208169 102 -208157
rect -46 -208207 46 -208201
rect -46 -208241 -34 -208207
rect 34 -208241 46 -208207
rect -46 -208247 46 -208241
rect -46 -208315 46 -208309
rect -46 -208349 -34 -208315
rect 34 -208349 46 -208315
rect -46 -208355 46 -208349
rect -102 -208399 -56 -208387
rect -102 -209375 -96 -208399
rect -62 -209375 -56 -208399
rect -102 -209387 -56 -209375
rect 56 -208399 102 -208387
rect 56 -209375 62 -208399
rect 96 -209375 102 -208399
rect 56 -209387 102 -209375
rect -46 -209425 46 -209419
rect -46 -209459 -34 -209425
rect 34 -209459 46 -209425
rect -46 -209465 46 -209459
rect -46 -209533 46 -209527
rect -46 -209567 -34 -209533
rect 34 -209567 46 -209533
rect -46 -209573 46 -209567
rect -102 -209617 -56 -209605
rect -102 -210593 -96 -209617
rect -62 -210593 -56 -209617
rect -102 -210605 -56 -210593
rect 56 -209617 102 -209605
rect 56 -210593 62 -209617
rect 96 -210593 102 -209617
rect 56 -210605 102 -210593
rect -46 -210643 46 -210637
rect -46 -210677 -34 -210643
rect 34 -210677 46 -210643
rect -46 -210683 46 -210677
rect -46 -210751 46 -210745
rect -46 -210785 -34 -210751
rect 34 -210785 46 -210751
rect -46 -210791 46 -210785
rect -102 -210835 -56 -210823
rect -102 -211811 -96 -210835
rect -62 -211811 -56 -210835
rect -102 -211823 -56 -211811
rect 56 -210835 102 -210823
rect 56 -211811 62 -210835
rect 96 -211811 102 -210835
rect 56 -211823 102 -211811
rect -46 -211861 46 -211855
rect -46 -211895 -34 -211861
rect 34 -211895 46 -211861
rect -46 -211901 46 -211895
rect -46 -211969 46 -211963
rect -46 -212003 -34 -211969
rect 34 -212003 46 -211969
rect -46 -212009 46 -212003
rect -102 -212053 -56 -212041
rect -102 -213029 -96 -212053
rect -62 -213029 -56 -212053
rect -102 -213041 -56 -213029
rect 56 -212053 102 -212041
rect 56 -213029 62 -212053
rect 96 -213029 102 -212053
rect 56 -213041 102 -213029
rect -46 -213079 46 -213073
rect -46 -213113 -34 -213079
rect 34 -213113 46 -213079
rect -46 -213119 46 -213113
rect -46 -213187 46 -213181
rect -46 -213221 -34 -213187
rect 34 -213221 46 -213187
rect -46 -213227 46 -213221
rect -102 -213271 -56 -213259
rect -102 -214247 -96 -213271
rect -62 -214247 -56 -213271
rect -102 -214259 -56 -214247
rect 56 -213271 102 -213259
rect 56 -214247 62 -213271
rect 96 -214247 102 -213271
rect 56 -214259 102 -214247
rect -46 -214297 46 -214291
rect -46 -214331 -34 -214297
rect 34 -214331 46 -214297
rect -46 -214337 46 -214331
rect -46 -214405 46 -214399
rect -46 -214439 -34 -214405
rect 34 -214439 46 -214405
rect -46 -214445 46 -214439
rect -102 -214489 -56 -214477
rect -102 -215465 -96 -214489
rect -62 -215465 -56 -214489
rect -102 -215477 -56 -215465
rect 56 -214489 102 -214477
rect 56 -215465 62 -214489
rect 96 -215465 102 -214489
rect 56 -215477 102 -215465
rect -46 -215515 46 -215509
rect -46 -215549 -34 -215515
rect 34 -215549 46 -215515
rect -46 -215555 46 -215549
rect -46 -215623 46 -215617
rect -46 -215657 -34 -215623
rect 34 -215657 46 -215623
rect -46 -215663 46 -215657
rect -102 -215707 -56 -215695
rect -102 -216683 -96 -215707
rect -62 -216683 -56 -215707
rect -102 -216695 -56 -216683
rect 56 -215707 102 -215695
rect 56 -216683 62 -215707
rect 96 -216683 102 -215707
rect 56 -216695 102 -216683
rect -46 -216733 46 -216727
rect -46 -216767 -34 -216733
rect 34 -216767 46 -216733
rect -46 -216773 46 -216767
rect -46 -216841 46 -216835
rect -46 -216875 -34 -216841
rect 34 -216875 46 -216841
rect -46 -216881 46 -216875
rect -102 -216925 -56 -216913
rect -102 -217901 -96 -216925
rect -62 -217901 -56 -216925
rect -102 -217913 -56 -217901
rect 56 -216925 102 -216913
rect 56 -217901 62 -216925
rect 96 -217901 102 -216925
rect 56 -217913 102 -217901
rect -46 -217951 46 -217945
rect -46 -217985 -34 -217951
rect 34 -217985 46 -217951
rect -46 -217991 46 -217985
rect -46 -218059 46 -218053
rect -46 -218093 -34 -218059
rect 34 -218093 46 -218059
rect -46 -218099 46 -218093
rect -102 -218143 -56 -218131
rect -102 -219119 -96 -218143
rect -62 -219119 -56 -218143
rect -102 -219131 -56 -219119
rect 56 -218143 102 -218131
rect 56 -219119 62 -218143
rect 96 -219119 102 -218143
rect 56 -219131 102 -219119
rect -46 -219169 46 -219163
rect -46 -219203 -34 -219169
rect 34 -219203 46 -219169
rect -46 -219209 46 -219203
rect -46 -219277 46 -219271
rect -46 -219311 -34 -219277
rect 34 -219311 46 -219277
rect -46 -219317 46 -219311
rect -102 -219361 -56 -219349
rect -102 -220337 -96 -219361
rect -62 -220337 -56 -219361
rect -102 -220349 -56 -220337
rect 56 -219361 102 -219349
rect 56 -220337 62 -219361
rect 96 -220337 102 -219361
rect 56 -220349 102 -220337
rect -46 -220387 46 -220381
rect -46 -220421 -34 -220387
rect 34 -220421 46 -220387
rect -46 -220427 46 -220421
rect -46 -220495 46 -220489
rect -46 -220529 -34 -220495
rect 34 -220529 46 -220495
rect -46 -220535 46 -220529
rect -102 -220579 -56 -220567
rect -102 -221555 -96 -220579
rect -62 -221555 -56 -220579
rect -102 -221567 -56 -221555
rect 56 -220579 102 -220567
rect 56 -221555 62 -220579
rect 96 -221555 102 -220579
rect 56 -221567 102 -221555
rect -46 -221605 46 -221599
rect -46 -221639 -34 -221605
rect 34 -221639 46 -221605
rect -46 -221645 46 -221639
rect -46 -221713 46 -221707
rect -46 -221747 -34 -221713
rect 34 -221747 46 -221713
rect -46 -221753 46 -221747
rect -102 -221797 -56 -221785
rect -102 -222773 -96 -221797
rect -62 -222773 -56 -221797
rect -102 -222785 -56 -222773
rect 56 -221797 102 -221785
rect 56 -222773 62 -221797
rect 96 -222773 102 -221797
rect 56 -222785 102 -222773
rect -46 -222823 46 -222817
rect -46 -222857 -34 -222823
rect 34 -222857 46 -222823
rect -46 -222863 46 -222857
rect -46 -222931 46 -222925
rect -46 -222965 -34 -222931
rect 34 -222965 46 -222931
rect -46 -222971 46 -222965
rect -102 -223015 -56 -223003
rect -102 -223991 -96 -223015
rect -62 -223991 -56 -223015
rect -102 -224003 -56 -223991
rect 56 -223015 102 -223003
rect 56 -223991 62 -223015
rect 96 -223991 102 -223015
rect 56 -224003 102 -223991
rect -46 -224041 46 -224035
rect -46 -224075 -34 -224041
rect 34 -224075 46 -224041
rect -46 -224081 46 -224075
rect -46 -224149 46 -224143
rect -46 -224183 -34 -224149
rect 34 -224183 46 -224149
rect -46 -224189 46 -224183
rect -102 -224233 -56 -224221
rect -102 -225209 -96 -224233
rect -62 -225209 -56 -224233
rect -102 -225221 -56 -225209
rect 56 -224233 102 -224221
rect 56 -225209 62 -224233
rect 96 -225209 102 -224233
rect 56 -225221 102 -225209
rect -46 -225259 46 -225253
rect -46 -225293 -34 -225259
rect 34 -225293 46 -225259
rect -46 -225299 46 -225293
rect -46 -225367 46 -225361
rect -46 -225401 -34 -225367
rect 34 -225401 46 -225367
rect -46 -225407 46 -225401
rect -102 -225451 -56 -225439
rect -102 -226427 -96 -225451
rect -62 -226427 -56 -225451
rect -102 -226439 -56 -226427
rect 56 -225451 102 -225439
rect 56 -226427 62 -225451
rect 96 -226427 102 -225451
rect 56 -226439 102 -226427
rect -46 -226477 46 -226471
rect -46 -226511 -34 -226477
rect 34 -226511 46 -226477
rect -46 -226517 46 -226511
rect -46 -226585 46 -226579
rect -46 -226619 -34 -226585
rect 34 -226619 46 -226585
rect -46 -226625 46 -226619
rect -102 -226669 -56 -226657
rect -102 -227645 -96 -226669
rect -62 -227645 -56 -226669
rect -102 -227657 -56 -227645
rect 56 -226669 102 -226657
rect 56 -227645 62 -226669
rect 96 -227645 102 -226669
rect 56 -227657 102 -227645
rect -46 -227695 46 -227689
rect -46 -227729 -34 -227695
rect 34 -227729 46 -227695
rect -46 -227735 46 -227729
rect -46 -227803 46 -227797
rect -46 -227837 -34 -227803
rect 34 -227837 46 -227803
rect -46 -227843 46 -227837
rect -102 -227887 -56 -227875
rect -102 -228863 -96 -227887
rect -62 -228863 -56 -227887
rect -102 -228875 -56 -228863
rect 56 -227887 102 -227875
rect 56 -228863 62 -227887
rect 96 -228863 102 -227887
rect 56 -228875 102 -228863
rect -46 -228913 46 -228907
rect -46 -228947 -34 -228913
rect 34 -228947 46 -228913
rect -46 -228953 46 -228947
rect -46 -229021 46 -229015
rect -46 -229055 -34 -229021
rect 34 -229055 46 -229021
rect -46 -229061 46 -229055
rect -102 -229105 -56 -229093
rect -102 -230081 -96 -229105
rect -62 -230081 -56 -229105
rect -102 -230093 -56 -230081
rect 56 -229105 102 -229093
rect 56 -230081 62 -229105
rect 96 -230081 102 -229105
rect 56 -230093 102 -230081
rect -46 -230131 46 -230125
rect -46 -230165 -34 -230131
rect 34 -230165 46 -230131
rect -46 -230171 46 -230165
rect -46 -230239 46 -230233
rect -46 -230273 -34 -230239
rect 34 -230273 46 -230239
rect -46 -230279 46 -230273
rect -102 -230323 -56 -230311
rect -102 -231299 -96 -230323
rect -62 -231299 -56 -230323
rect -102 -231311 -56 -231299
rect 56 -230323 102 -230311
rect 56 -231299 62 -230323
rect 96 -231299 102 -230323
rect 56 -231311 102 -231299
rect -46 -231349 46 -231343
rect -46 -231383 -34 -231349
rect 34 -231383 46 -231349
rect -46 -231389 46 -231383
rect -46 -231457 46 -231451
rect -46 -231491 -34 -231457
rect 34 -231491 46 -231457
rect -46 -231497 46 -231491
rect -102 -231541 -56 -231529
rect -102 -232517 -96 -231541
rect -62 -232517 -56 -231541
rect -102 -232529 -56 -232517
rect 56 -231541 102 -231529
rect 56 -232517 62 -231541
rect 96 -232517 102 -231541
rect 56 -232529 102 -232517
rect -46 -232567 46 -232561
rect -46 -232601 -34 -232567
rect 34 -232601 46 -232567
rect -46 -232607 46 -232601
rect -46 -232675 46 -232669
rect -46 -232709 -34 -232675
rect 34 -232709 46 -232675
rect -46 -232715 46 -232709
rect -102 -232759 -56 -232747
rect -102 -233735 -96 -232759
rect -62 -233735 -56 -232759
rect -102 -233747 -56 -233735
rect 56 -232759 102 -232747
rect 56 -233735 62 -232759
rect 96 -233735 102 -232759
rect 56 -233747 102 -233735
rect -46 -233785 46 -233779
rect -46 -233819 -34 -233785
rect 34 -233819 46 -233785
rect -46 -233825 46 -233819
rect -46 -233893 46 -233887
rect -46 -233927 -34 -233893
rect 34 -233927 46 -233893
rect -46 -233933 46 -233927
rect -102 -233977 -56 -233965
rect -102 -234953 -96 -233977
rect -62 -234953 -56 -233977
rect -102 -234965 -56 -234953
rect 56 -233977 102 -233965
rect 56 -234953 62 -233977
rect 96 -234953 102 -233977
rect 56 -234965 102 -234953
rect -46 -235003 46 -234997
rect -46 -235037 -34 -235003
rect 34 -235037 46 -235003
rect -46 -235043 46 -235037
rect -46 -235111 46 -235105
rect -46 -235145 -34 -235111
rect 34 -235145 46 -235111
rect -46 -235151 46 -235145
rect -102 -235195 -56 -235183
rect -102 -236171 -96 -235195
rect -62 -236171 -56 -235195
rect -102 -236183 -56 -236171
rect 56 -235195 102 -235183
rect 56 -236171 62 -235195
rect 96 -236171 102 -235195
rect 56 -236183 102 -236171
rect -46 -236221 46 -236215
rect -46 -236255 -34 -236221
rect 34 -236255 46 -236221
rect -46 -236261 46 -236255
rect -46 -236329 46 -236323
rect -46 -236363 -34 -236329
rect 34 -236363 46 -236329
rect -46 -236369 46 -236363
rect -102 -236413 -56 -236401
rect -102 -237389 -96 -236413
rect -62 -237389 -56 -236413
rect -102 -237401 -56 -237389
rect 56 -236413 102 -236401
rect 56 -237389 62 -236413
rect 96 -237389 102 -236413
rect 56 -237401 102 -237389
rect -46 -237439 46 -237433
rect -46 -237473 -34 -237439
rect 34 -237473 46 -237439
rect -46 -237479 46 -237473
rect -46 -237547 46 -237541
rect -46 -237581 -34 -237547
rect 34 -237581 46 -237547
rect -46 -237587 46 -237581
rect -102 -237631 -56 -237619
rect -102 -238607 -96 -237631
rect -62 -238607 -56 -237631
rect -102 -238619 -56 -238607
rect 56 -237631 102 -237619
rect 56 -238607 62 -237631
rect 96 -238607 102 -237631
rect 56 -238619 102 -238607
rect -46 -238657 46 -238651
rect -46 -238691 -34 -238657
rect 34 -238691 46 -238657
rect -46 -238697 46 -238691
rect -46 -238765 46 -238759
rect -46 -238799 -34 -238765
rect 34 -238799 46 -238765
rect -46 -238805 46 -238799
rect -102 -238849 -56 -238837
rect -102 -239825 -96 -238849
rect -62 -239825 -56 -238849
rect -102 -239837 -56 -239825
rect 56 -238849 102 -238837
rect 56 -239825 62 -238849
rect 96 -239825 102 -238849
rect 56 -239837 102 -239825
rect -46 -239875 46 -239869
rect -46 -239909 -34 -239875
rect 34 -239909 46 -239875
rect -46 -239915 46 -239909
rect -46 -239983 46 -239977
rect -46 -240017 -34 -239983
rect 34 -240017 46 -239983
rect -46 -240023 46 -240017
rect -102 -240067 -56 -240055
rect -102 -241043 -96 -240067
rect -62 -241043 -56 -240067
rect -102 -241055 -56 -241043
rect 56 -240067 102 -240055
rect 56 -241043 62 -240067
rect 96 -241043 102 -240067
rect 56 -241055 102 -241043
rect -46 -241093 46 -241087
rect -46 -241127 -34 -241093
rect 34 -241127 46 -241093
rect -46 -241133 46 -241127
rect -46 -241201 46 -241195
rect -46 -241235 -34 -241201
rect 34 -241235 46 -241201
rect -46 -241241 46 -241235
rect -102 -241285 -56 -241273
rect -102 -242261 -96 -241285
rect -62 -242261 -56 -241285
rect -102 -242273 -56 -242261
rect 56 -241285 102 -241273
rect 56 -242261 62 -241285
rect 96 -242261 102 -241285
rect 56 -242273 102 -242261
rect -46 -242311 46 -242305
rect -46 -242345 -34 -242311
rect 34 -242345 46 -242311
rect -46 -242351 46 -242345
rect -46 -242419 46 -242413
rect -46 -242453 -34 -242419
rect 34 -242453 46 -242419
rect -46 -242459 46 -242453
rect -102 -242503 -56 -242491
rect -102 -243479 -96 -242503
rect -62 -243479 -56 -242503
rect -102 -243491 -56 -243479
rect 56 -242503 102 -242491
rect 56 -243479 62 -242503
rect 96 -243479 102 -242503
rect 56 -243491 102 -243479
rect -46 -243529 46 -243523
rect -46 -243563 -34 -243529
rect 34 -243563 46 -243529
rect -46 -243569 46 -243563
rect -46 -243637 46 -243631
rect -46 -243671 -34 -243637
rect 34 -243671 46 -243637
rect -46 -243677 46 -243671
rect -102 -243721 -56 -243709
rect -102 -244697 -96 -243721
rect -62 -244697 -56 -243721
rect -102 -244709 -56 -244697
rect 56 -243721 102 -243709
rect 56 -244697 62 -243721
rect 96 -244697 102 -243721
rect 56 -244709 102 -244697
rect -46 -244747 46 -244741
rect -46 -244781 -34 -244747
rect 34 -244781 46 -244747
rect -46 -244787 46 -244781
rect -46 -244855 46 -244849
rect -46 -244889 -34 -244855
rect 34 -244889 46 -244855
rect -46 -244895 46 -244889
rect -102 -244939 -56 -244927
rect -102 -245915 -96 -244939
rect -62 -245915 -56 -244939
rect -102 -245927 -56 -245915
rect 56 -244939 102 -244927
rect 56 -245915 62 -244939
rect 96 -245915 102 -244939
rect 56 -245927 102 -245915
rect -46 -245965 46 -245959
rect -46 -245999 -34 -245965
rect 34 -245999 46 -245965
rect -46 -246005 46 -245999
rect -46 -246073 46 -246067
rect -46 -246107 -34 -246073
rect 34 -246107 46 -246073
rect -46 -246113 46 -246107
rect -102 -246157 -56 -246145
rect -102 -247133 -96 -246157
rect -62 -247133 -56 -246157
rect -102 -247145 -56 -247133
rect 56 -246157 102 -246145
rect 56 -247133 62 -246157
rect 96 -247133 102 -246157
rect 56 -247145 102 -247133
rect -46 -247183 46 -247177
rect -46 -247217 -34 -247183
rect 34 -247217 46 -247183
rect -46 -247223 46 -247217
rect -46 -247291 46 -247285
rect -46 -247325 -34 -247291
rect 34 -247325 46 -247291
rect -46 -247331 46 -247325
rect -102 -247375 -56 -247363
rect -102 -248351 -96 -247375
rect -62 -248351 -56 -247375
rect -102 -248363 -56 -248351
rect 56 -247375 102 -247363
rect 56 -248351 62 -247375
rect 96 -248351 102 -247375
rect 56 -248363 102 -248351
rect -46 -248401 46 -248395
rect -46 -248435 -34 -248401
rect 34 -248435 46 -248401
rect -46 -248441 46 -248435
rect -46 -248509 46 -248503
rect -46 -248543 -34 -248509
rect 34 -248543 46 -248509
rect -46 -248549 46 -248543
rect -102 -248593 -56 -248581
rect -102 -249569 -96 -248593
rect -62 -249569 -56 -248593
rect -102 -249581 -56 -249569
rect 56 -248593 102 -248581
rect 56 -249569 62 -248593
rect 96 -249569 102 -248593
rect 56 -249581 102 -249569
rect -46 -249619 46 -249613
rect -46 -249653 -34 -249619
rect 34 -249653 46 -249619
rect -46 -249659 46 -249653
rect -46 -249727 46 -249721
rect -46 -249761 -34 -249727
rect 34 -249761 46 -249727
rect -46 -249767 46 -249761
rect -102 -249811 -56 -249799
rect -102 -250787 -96 -249811
rect -62 -250787 -56 -249811
rect -102 -250799 -56 -250787
rect 56 -249811 102 -249799
rect 56 -250787 62 -249811
rect 96 -250787 102 -249811
rect 56 -250799 102 -250787
rect -46 -250837 46 -250831
rect -46 -250871 -34 -250837
rect 34 -250871 46 -250837
rect -46 -250877 46 -250871
rect -46 -250945 46 -250939
rect -46 -250979 -34 -250945
rect 34 -250979 46 -250945
rect -46 -250985 46 -250979
rect -102 -251029 -56 -251017
rect -102 -252005 -96 -251029
rect -62 -252005 -56 -251029
rect -102 -252017 -56 -252005
rect 56 -251029 102 -251017
rect 56 -252005 62 -251029
rect 96 -252005 102 -251029
rect 56 -252017 102 -252005
rect -46 -252055 46 -252049
rect -46 -252089 -34 -252055
rect 34 -252089 46 -252055
rect -46 -252095 46 -252089
rect -46 -252163 46 -252157
rect -46 -252197 -34 -252163
rect 34 -252197 46 -252163
rect -46 -252203 46 -252197
rect -102 -252247 -56 -252235
rect -102 -253223 -96 -252247
rect -62 -253223 -56 -252247
rect -102 -253235 -56 -253223
rect 56 -252247 102 -252235
rect 56 -253223 62 -252247
rect 96 -253223 102 -252247
rect 56 -253235 102 -253223
rect -46 -253273 46 -253267
rect -46 -253307 -34 -253273
rect 34 -253307 46 -253273
rect -46 -253313 46 -253307
rect -46 -253381 46 -253375
rect -46 -253415 -34 -253381
rect 34 -253415 46 -253381
rect -46 -253421 46 -253415
rect -102 -253465 -56 -253453
rect -102 -254441 -96 -253465
rect -62 -254441 -56 -253465
rect -102 -254453 -56 -254441
rect 56 -253465 102 -253453
rect 56 -254441 62 -253465
rect 96 -254441 102 -253465
rect 56 -254453 102 -254441
rect -46 -254491 46 -254485
rect -46 -254525 -34 -254491
rect 34 -254525 46 -254491
rect -46 -254531 46 -254525
rect -46 -254599 46 -254593
rect -46 -254633 -34 -254599
rect 34 -254633 46 -254599
rect -46 -254639 46 -254633
rect -102 -254683 -56 -254671
rect -102 -255659 -96 -254683
rect -62 -255659 -56 -254683
rect -102 -255671 -56 -255659
rect 56 -254683 102 -254671
rect 56 -255659 62 -254683
rect 96 -255659 102 -254683
rect 56 -255671 102 -255659
rect -46 -255709 46 -255703
rect -46 -255743 -34 -255709
rect 34 -255743 46 -255709
rect -46 -255749 46 -255743
rect -46 -255817 46 -255811
rect -46 -255851 -34 -255817
rect 34 -255851 46 -255817
rect -46 -255857 46 -255851
rect -102 -255901 -56 -255889
rect -102 -256877 -96 -255901
rect -62 -256877 -56 -255901
rect -102 -256889 -56 -256877
rect 56 -255901 102 -255889
rect 56 -256877 62 -255901
rect 96 -256877 102 -255901
rect 56 -256889 102 -256877
rect -46 -256927 46 -256921
rect -46 -256961 -34 -256927
rect 34 -256961 46 -256927
rect -46 -256967 46 -256961
rect -46 -257035 46 -257029
rect -46 -257069 -34 -257035
rect 34 -257069 46 -257035
rect -46 -257075 46 -257069
rect -102 -257119 -56 -257107
rect -102 -258095 -96 -257119
rect -62 -258095 -56 -257119
rect -102 -258107 -56 -258095
rect 56 -257119 102 -257107
rect 56 -258095 62 -257119
rect 96 -258095 102 -257119
rect 56 -258107 102 -258095
rect -46 -258145 46 -258139
rect -46 -258179 -34 -258145
rect 34 -258179 46 -258145
rect -46 -258185 46 -258179
rect -46 -258253 46 -258247
rect -46 -258287 -34 -258253
rect 34 -258287 46 -258253
rect -46 -258293 46 -258287
rect -102 -258337 -56 -258325
rect -102 -259313 -96 -258337
rect -62 -259313 -56 -258337
rect -102 -259325 -56 -259313
rect 56 -258337 102 -258325
rect 56 -259313 62 -258337
rect 96 -259313 102 -258337
rect 56 -259325 102 -259313
rect -46 -259363 46 -259357
rect -46 -259397 -34 -259363
rect 34 -259397 46 -259363
rect -46 -259403 46 -259397
rect -46 -259471 46 -259465
rect -46 -259505 -34 -259471
rect 34 -259505 46 -259471
rect -46 -259511 46 -259505
rect -102 -259555 -56 -259543
rect -102 -260531 -96 -259555
rect -62 -260531 -56 -259555
rect -102 -260543 -56 -260531
rect 56 -259555 102 -259543
rect 56 -260531 62 -259555
rect 96 -260531 102 -259555
rect 56 -260543 102 -260531
rect -46 -260581 46 -260575
rect -46 -260615 -34 -260581
rect 34 -260615 46 -260581
rect -46 -260621 46 -260615
rect -46 -260689 46 -260683
rect -46 -260723 -34 -260689
rect 34 -260723 46 -260689
rect -46 -260729 46 -260723
rect -102 -260773 -56 -260761
rect -102 -261749 -96 -260773
rect -62 -261749 -56 -260773
rect -102 -261761 -56 -261749
rect 56 -260773 102 -260761
rect 56 -261749 62 -260773
rect 96 -261749 102 -260773
rect 56 -261761 102 -261749
rect -46 -261799 46 -261793
rect -46 -261833 -34 -261799
rect 34 -261833 46 -261799
rect -46 -261839 46 -261833
rect -46 -261907 46 -261901
rect -46 -261941 -34 -261907
rect 34 -261941 46 -261907
rect -46 -261947 46 -261941
rect -102 -261991 -56 -261979
rect -102 -262967 -96 -261991
rect -62 -262967 -56 -261991
rect -102 -262979 -56 -262967
rect 56 -261991 102 -261979
rect 56 -262967 62 -261991
rect 96 -262967 102 -261991
rect 56 -262979 102 -262967
rect -46 -263017 46 -263011
rect -46 -263051 -34 -263017
rect 34 -263051 46 -263017
rect -46 -263057 46 -263051
rect -46 -263125 46 -263119
rect -46 -263159 -34 -263125
rect 34 -263159 46 -263125
rect -46 -263165 46 -263159
rect -102 -263209 -56 -263197
rect -102 -264185 -96 -263209
rect -62 -264185 -56 -263209
rect -102 -264197 -56 -264185
rect 56 -263209 102 -263197
rect 56 -264185 62 -263209
rect 96 -264185 102 -263209
rect 56 -264197 102 -264185
rect -46 -264235 46 -264229
rect -46 -264269 -34 -264235
rect 34 -264269 46 -264235
rect -46 -264275 46 -264269
rect -46 -264343 46 -264337
rect -46 -264377 -34 -264343
rect 34 -264377 46 -264343
rect -46 -264383 46 -264377
rect -102 -264427 -56 -264415
rect -102 -265403 -96 -264427
rect -62 -265403 -56 -264427
rect -102 -265415 -56 -265403
rect 56 -264427 102 -264415
rect 56 -265403 62 -264427
rect 96 -265403 102 -264427
rect 56 -265415 102 -265403
rect -46 -265453 46 -265447
rect -46 -265487 -34 -265453
rect 34 -265487 46 -265453
rect -46 -265493 46 -265487
rect -46 -265561 46 -265555
rect -46 -265595 -34 -265561
rect 34 -265595 46 -265561
rect -46 -265601 46 -265595
rect -102 -265645 -56 -265633
rect -102 -266621 -96 -265645
rect -62 -266621 -56 -265645
rect -102 -266633 -56 -266621
rect 56 -265645 102 -265633
rect 56 -266621 62 -265645
rect 96 -266621 102 -265645
rect 56 -266633 102 -266621
rect -46 -266671 46 -266665
rect -46 -266705 -34 -266671
rect 34 -266705 46 -266671
rect -46 -266711 46 -266705
rect -46 -266779 46 -266773
rect -46 -266813 -34 -266779
rect 34 -266813 46 -266779
rect -46 -266819 46 -266813
rect -102 -266863 -56 -266851
rect -102 -267839 -96 -266863
rect -62 -267839 -56 -266863
rect -102 -267851 -56 -267839
rect 56 -266863 102 -266851
rect 56 -267839 62 -266863
rect 96 -267839 102 -266863
rect 56 -267851 102 -267839
rect -46 -267889 46 -267883
rect -46 -267923 -34 -267889
rect 34 -267923 46 -267889
rect -46 -267929 46 -267923
rect -46 -267997 46 -267991
rect -46 -268031 -34 -267997
rect 34 -268031 46 -267997
rect -46 -268037 46 -268031
rect -102 -268081 -56 -268069
rect -102 -269057 -96 -268081
rect -62 -269057 -56 -268081
rect -102 -269069 -56 -269057
rect 56 -268081 102 -268069
rect 56 -269057 62 -268081
rect 96 -269057 102 -268081
rect 56 -269069 102 -269057
rect -46 -269107 46 -269101
rect -46 -269141 -34 -269107
rect 34 -269141 46 -269107
rect -46 -269147 46 -269141
rect -46 -269215 46 -269209
rect -46 -269249 -34 -269215
rect 34 -269249 46 -269215
rect -46 -269255 46 -269249
rect -102 -269299 -56 -269287
rect -102 -270275 -96 -269299
rect -62 -270275 -56 -269299
rect -102 -270287 -56 -270275
rect 56 -269299 102 -269287
rect 56 -270275 62 -269299
rect 96 -270275 102 -269299
rect 56 -270287 102 -270275
rect -46 -270325 46 -270319
rect -46 -270359 -34 -270325
rect 34 -270359 46 -270325
rect -46 -270365 46 -270359
rect -46 -270433 46 -270427
rect -46 -270467 -34 -270433
rect 34 -270467 46 -270433
rect -46 -270473 46 -270467
rect -102 -270517 -56 -270505
rect -102 -271493 -96 -270517
rect -62 -271493 -56 -270517
rect -102 -271505 -56 -271493
rect 56 -270517 102 -270505
rect 56 -271493 62 -270517
rect 96 -271493 102 -270517
rect 56 -271505 102 -271493
rect -46 -271543 46 -271537
rect -46 -271577 -34 -271543
rect 34 -271577 46 -271543
rect -46 -271583 46 -271577
rect -46 -271651 46 -271645
rect -46 -271685 -34 -271651
rect 34 -271685 46 -271651
rect -46 -271691 46 -271685
rect -102 -271735 -56 -271723
rect -102 -272711 -96 -271735
rect -62 -272711 -56 -271735
rect -102 -272723 -56 -272711
rect 56 -271735 102 -271723
rect 56 -272711 62 -271735
rect 96 -272711 102 -271735
rect 56 -272723 102 -272711
rect -46 -272761 46 -272755
rect -46 -272795 -34 -272761
rect 34 -272795 46 -272761
rect -46 -272801 46 -272795
rect -46 -272869 46 -272863
rect -46 -272903 -34 -272869
rect 34 -272903 46 -272869
rect -46 -272909 46 -272903
rect -102 -272953 -56 -272941
rect -102 -273929 -96 -272953
rect -62 -273929 -56 -272953
rect -102 -273941 -56 -273929
rect 56 -272953 102 -272941
rect 56 -273929 62 -272953
rect 96 -273929 102 -272953
rect 56 -273941 102 -273929
rect -46 -273979 46 -273973
rect -46 -274013 -34 -273979
rect 34 -274013 46 -273979
rect -46 -274019 46 -274013
rect -46 -274087 46 -274081
rect -46 -274121 -34 -274087
rect 34 -274121 46 -274087
rect -46 -274127 46 -274121
rect -102 -274171 -56 -274159
rect -102 -275147 -96 -274171
rect -62 -275147 -56 -274171
rect -102 -275159 -56 -275147
rect 56 -274171 102 -274159
rect 56 -275147 62 -274171
rect 96 -275147 102 -274171
rect 56 -275159 102 -275147
rect -46 -275197 46 -275191
rect -46 -275231 -34 -275197
rect 34 -275231 46 -275197
rect -46 -275237 46 -275231
rect -46 -275305 46 -275299
rect -46 -275339 -34 -275305
rect 34 -275339 46 -275305
rect -46 -275345 46 -275339
rect -102 -275389 -56 -275377
rect -102 -276365 -96 -275389
rect -62 -276365 -56 -275389
rect -102 -276377 -56 -276365
rect 56 -275389 102 -275377
rect 56 -276365 62 -275389
rect 96 -276365 102 -275389
rect 56 -276377 102 -276365
rect -46 -276415 46 -276409
rect -46 -276449 -34 -276415
rect 34 -276449 46 -276415
rect -46 -276455 46 -276449
rect -46 -276523 46 -276517
rect -46 -276557 -34 -276523
rect 34 -276557 46 -276523
rect -46 -276563 46 -276557
rect -102 -276607 -56 -276595
rect -102 -277583 -96 -276607
rect -62 -277583 -56 -276607
rect -102 -277595 -56 -277583
rect 56 -276607 102 -276595
rect 56 -277583 62 -276607
rect 96 -277583 102 -276607
rect 56 -277595 102 -277583
rect -46 -277633 46 -277627
rect -46 -277667 -34 -277633
rect 34 -277667 46 -277633
rect -46 -277673 46 -277667
rect -46 -277741 46 -277735
rect -46 -277775 -34 -277741
rect 34 -277775 46 -277741
rect -46 -277781 46 -277775
rect -102 -277825 -56 -277813
rect -102 -278801 -96 -277825
rect -62 -278801 -56 -277825
rect -102 -278813 -56 -278801
rect 56 -277825 102 -277813
rect 56 -278801 62 -277825
rect 96 -278801 102 -277825
rect 56 -278813 102 -278801
rect -46 -278851 46 -278845
rect -46 -278885 -34 -278851
rect 34 -278885 46 -278851
rect -46 -278891 46 -278885
rect -46 -278959 46 -278953
rect -46 -278993 -34 -278959
rect 34 -278993 46 -278959
rect -46 -278999 46 -278993
rect -102 -279043 -56 -279031
rect -102 -280019 -96 -279043
rect -62 -280019 -56 -279043
rect -102 -280031 -56 -280019
rect 56 -279043 102 -279031
rect 56 -280019 62 -279043
rect 96 -280019 102 -279043
rect 56 -280031 102 -280019
rect -46 -280069 46 -280063
rect -46 -280103 -34 -280069
rect 34 -280103 46 -280069
rect -46 -280109 46 -280103
rect -46 -280177 46 -280171
rect -46 -280211 -34 -280177
rect 34 -280211 46 -280177
rect -46 -280217 46 -280211
rect -102 -280261 -56 -280249
rect -102 -281237 -96 -280261
rect -62 -281237 -56 -280261
rect -102 -281249 -56 -281237
rect 56 -280261 102 -280249
rect 56 -281237 62 -280261
rect 96 -281237 102 -280261
rect 56 -281249 102 -281237
rect -46 -281287 46 -281281
rect -46 -281321 -34 -281287
rect 34 -281321 46 -281287
rect -46 -281327 46 -281321
rect -46 -281395 46 -281389
rect -46 -281429 -34 -281395
rect 34 -281429 46 -281395
rect -46 -281435 46 -281429
rect -102 -281479 -56 -281467
rect -102 -282455 -96 -281479
rect -62 -282455 -56 -281479
rect -102 -282467 -56 -282455
rect 56 -281479 102 -281467
rect 56 -282455 62 -281479
rect 96 -282455 102 -281479
rect 56 -282467 102 -282455
rect -46 -282505 46 -282499
rect -46 -282539 -34 -282505
rect 34 -282539 46 -282505
rect -46 -282545 46 -282539
rect -46 -282613 46 -282607
rect -46 -282647 -34 -282613
rect 34 -282647 46 -282613
rect -46 -282653 46 -282647
rect -102 -282697 -56 -282685
rect -102 -283673 -96 -282697
rect -62 -283673 -56 -282697
rect -102 -283685 -56 -283673
rect 56 -282697 102 -282685
rect 56 -283673 62 -282697
rect 96 -283673 102 -282697
rect 56 -283685 102 -283673
rect -46 -283723 46 -283717
rect -46 -283757 -34 -283723
rect 34 -283757 46 -283723
rect -46 -283763 46 -283757
rect -46 -283831 46 -283825
rect -46 -283865 -34 -283831
rect 34 -283865 46 -283831
rect -46 -283871 46 -283865
rect -102 -283915 -56 -283903
rect -102 -284891 -96 -283915
rect -62 -284891 -56 -283915
rect -102 -284903 -56 -284891
rect 56 -283915 102 -283903
rect 56 -284891 62 -283915
rect 96 -284891 102 -283915
rect 56 -284903 102 -284891
rect -46 -284941 46 -284935
rect -46 -284975 -34 -284941
rect 34 -284975 46 -284941
rect -46 -284981 46 -284975
rect -46 -285049 46 -285043
rect -46 -285083 -34 -285049
rect 34 -285083 46 -285049
rect -46 -285089 46 -285083
rect -102 -285133 -56 -285121
rect -102 -286109 -96 -285133
rect -62 -286109 -56 -285133
rect -102 -286121 -56 -286109
rect 56 -285133 102 -285121
rect 56 -286109 62 -285133
rect 96 -286109 102 -285133
rect 56 -286121 102 -286109
rect -46 -286159 46 -286153
rect -46 -286193 -34 -286159
rect 34 -286193 46 -286159
rect -46 -286199 46 -286193
rect -46 -286267 46 -286261
rect -46 -286301 -34 -286267
rect 34 -286301 46 -286267
rect -46 -286307 46 -286301
rect -102 -286351 -56 -286339
rect -102 -287327 -96 -286351
rect -62 -287327 -56 -286351
rect -102 -287339 -56 -287327
rect 56 -286351 102 -286339
rect 56 -287327 62 -286351
rect 96 -287327 102 -286351
rect 56 -287339 102 -287327
rect -46 -287377 46 -287371
rect -46 -287411 -34 -287377
rect 34 -287411 46 -287377
rect -46 -287417 46 -287411
rect -46 -287485 46 -287479
rect -46 -287519 -34 -287485
rect 34 -287519 46 -287485
rect -46 -287525 46 -287519
rect -102 -287569 -56 -287557
rect -102 -288545 -96 -287569
rect -62 -288545 -56 -287569
rect -102 -288557 -56 -288545
rect 56 -287569 102 -287557
rect 56 -288545 62 -287569
rect 96 -288545 102 -287569
rect 56 -288557 102 -288545
rect -46 -288595 46 -288589
rect -46 -288629 -34 -288595
rect 34 -288629 46 -288595
rect -46 -288635 46 -288629
rect -46 -288703 46 -288697
rect -46 -288737 -34 -288703
rect 34 -288737 46 -288703
rect -46 -288743 46 -288737
rect -102 -288787 -56 -288775
rect -102 -289763 -96 -288787
rect -62 -289763 -56 -288787
rect -102 -289775 -56 -289763
rect 56 -288787 102 -288775
rect 56 -289763 62 -288787
rect 96 -289763 102 -288787
rect 56 -289775 102 -289763
rect -46 -289813 46 -289807
rect -46 -289847 -34 -289813
rect 34 -289847 46 -289813
rect -46 -289853 46 -289847
rect -46 -289921 46 -289915
rect -46 -289955 -34 -289921
rect 34 -289955 46 -289921
rect -46 -289961 46 -289955
rect -102 -290005 -56 -289993
rect -102 -290981 -96 -290005
rect -62 -290981 -56 -290005
rect -102 -290993 -56 -290981
rect 56 -290005 102 -289993
rect 56 -290981 62 -290005
rect 96 -290981 102 -290005
rect 56 -290993 102 -290981
rect -46 -291031 46 -291025
rect -46 -291065 -34 -291031
rect 34 -291065 46 -291031
rect -46 -291071 46 -291065
rect -46 -291139 46 -291133
rect -46 -291173 -34 -291139
rect 34 -291173 46 -291139
rect -46 -291179 46 -291173
rect -102 -291223 -56 -291211
rect -102 -292199 -96 -291223
rect -62 -292199 -56 -291223
rect -102 -292211 -56 -292199
rect 56 -291223 102 -291211
rect 56 -292199 62 -291223
rect 96 -292199 102 -291223
rect 56 -292211 102 -292199
rect -46 -292249 46 -292243
rect -46 -292283 -34 -292249
rect 34 -292283 46 -292249
rect -46 -292289 46 -292283
rect -46 -292357 46 -292351
rect -46 -292391 -34 -292357
rect 34 -292391 46 -292357
rect -46 -292397 46 -292391
rect -102 -292441 -56 -292429
rect -102 -293417 -96 -292441
rect -62 -293417 -56 -292441
rect -102 -293429 -56 -293417
rect 56 -292441 102 -292429
rect 56 -293417 62 -292441
rect 96 -293417 102 -292441
rect 56 -293429 102 -293417
rect -46 -293467 46 -293461
rect -46 -293501 -34 -293467
rect 34 -293501 46 -293467
rect -46 -293507 46 -293501
rect -46 -293575 46 -293569
rect -46 -293609 -34 -293575
rect 34 -293609 46 -293575
rect -46 -293615 46 -293609
rect -102 -293659 -56 -293647
rect -102 -294635 -96 -293659
rect -62 -294635 -56 -293659
rect -102 -294647 -56 -294635
rect 56 -293659 102 -293647
rect 56 -294635 62 -293659
rect 96 -294635 102 -293659
rect 56 -294647 102 -294635
rect -46 -294685 46 -294679
rect -46 -294719 -34 -294685
rect 34 -294719 46 -294685
rect -46 -294725 46 -294719
rect -46 -294793 46 -294787
rect -46 -294827 -34 -294793
rect 34 -294827 46 -294793
rect -46 -294833 46 -294827
rect -102 -294877 -56 -294865
rect -102 -295853 -96 -294877
rect -62 -295853 -56 -294877
rect -102 -295865 -56 -295853
rect 56 -294877 102 -294865
rect 56 -295853 62 -294877
rect 96 -295853 102 -294877
rect 56 -295865 102 -295853
rect -46 -295903 46 -295897
rect -46 -295937 -34 -295903
rect 34 -295937 46 -295903
rect -46 -295943 46 -295937
rect -46 -296011 46 -296005
rect -46 -296045 -34 -296011
rect 34 -296045 46 -296011
rect -46 -296051 46 -296045
rect -102 -296095 -56 -296083
rect -102 -297071 -96 -296095
rect -62 -297071 -56 -296095
rect -102 -297083 -56 -297071
rect 56 -296095 102 -296083
rect 56 -297071 62 -296095
rect 96 -297071 102 -296095
rect 56 -297083 102 -297071
rect -46 -297121 46 -297115
rect -46 -297155 -34 -297121
rect 34 -297155 46 -297121
rect -46 -297161 46 -297155
rect -46 -297229 46 -297223
rect -46 -297263 -34 -297229
rect 34 -297263 46 -297229
rect -46 -297269 46 -297263
rect -102 -297313 -56 -297301
rect -102 -298289 -96 -297313
rect -62 -298289 -56 -297313
rect -102 -298301 -56 -298289
rect 56 -297313 102 -297301
rect 56 -298289 62 -297313
rect 96 -298289 102 -297313
rect 56 -298301 102 -298289
rect -46 -298339 46 -298333
rect -46 -298373 -34 -298339
rect 34 -298373 46 -298339
rect -46 -298379 46 -298373
rect -46 -298447 46 -298441
rect -46 -298481 -34 -298447
rect 34 -298481 46 -298447
rect -46 -298487 46 -298481
rect -102 -298531 -56 -298519
rect -102 -299507 -96 -298531
rect -62 -299507 -56 -298531
rect -102 -299519 -56 -299507
rect 56 -298531 102 -298519
rect 56 -299507 62 -298531
rect 96 -299507 102 -298531
rect 56 -299519 102 -299507
rect -46 -299557 46 -299551
rect -46 -299591 -34 -299557
rect 34 -299591 46 -299557
rect -46 -299597 46 -299591
rect -46 -299665 46 -299659
rect -46 -299699 -34 -299665
rect 34 -299699 46 -299665
rect -46 -299705 46 -299699
rect -102 -299749 -56 -299737
rect -102 -300725 -96 -299749
rect -62 -300725 -56 -299749
rect -102 -300737 -56 -300725
rect 56 -299749 102 -299737
rect 56 -300725 62 -299749
rect 96 -300725 102 -299749
rect 56 -300737 102 -300725
rect -46 -300775 46 -300769
rect -46 -300809 -34 -300775
rect 34 -300809 46 -300775
rect -46 -300815 46 -300809
rect -46 -300883 46 -300877
rect -46 -300917 -34 -300883
rect 34 -300917 46 -300883
rect -46 -300923 46 -300917
rect -102 -300967 -56 -300955
rect -102 -301943 -96 -300967
rect -62 -301943 -56 -300967
rect -102 -301955 -56 -301943
rect 56 -300967 102 -300955
rect 56 -301943 62 -300967
rect 96 -301943 102 -300967
rect 56 -301955 102 -301943
rect -46 -301993 46 -301987
rect -46 -302027 -34 -301993
rect 34 -302027 46 -301993
rect -46 -302033 46 -302027
rect -46 -302101 46 -302095
rect -46 -302135 -34 -302101
rect 34 -302135 46 -302101
rect -46 -302141 46 -302135
rect -102 -302185 -56 -302173
rect -102 -303161 -96 -302185
rect -62 -303161 -56 -302185
rect -102 -303173 -56 -303161
rect 56 -302185 102 -302173
rect 56 -303161 62 -302185
rect 96 -303161 102 -302185
rect 56 -303173 102 -303161
rect -46 -303211 46 -303205
rect -46 -303245 -34 -303211
rect 34 -303245 46 -303211
rect -46 -303251 46 -303245
rect -46 -303319 46 -303313
rect -46 -303353 -34 -303319
rect 34 -303353 46 -303319
rect -46 -303359 46 -303353
rect -102 -303403 -56 -303391
rect -102 -304379 -96 -303403
rect -62 -304379 -56 -303403
rect -102 -304391 -56 -304379
rect 56 -303403 102 -303391
rect 56 -304379 62 -303403
rect 96 -304379 102 -303403
rect 56 -304391 102 -304379
rect -46 -304429 46 -304423
rect -46 -304463 -34 -304429
rect 34 -304463 46 -304429
rect -46 -304469 46 -304463
rect -46 -304537 46 -304531
rect -46 -304571 -34 -304537
rect 34 -304571 46 -304537
rect -46 -304577 46 -304571
rect -102 -304621 -56 -304609
rect -102 -305597 -96 -304621
rect -62 -305597 -56 -304621
rect -102 -305609 -56 -305597
rect 56 -304621 102 -304609
rect 56 -305597 62 -304621
rect 96 -305597 102 -304621
rect 56 -305609 102 -305597
rect -46 -305647 46 -305641
rect -46 -305681 -34 -305647
rect 34 -305681 46 -305647
rect -46 -305687 46 -305681
rect -46 -305755 46 -305749
rect -46 -305789 -34 -305755
rect 34 -305789 46 -305755
rect -46 -305795 46 -305789
rect -102 -305839 -56 -305827
rect -102 -306815 -96 -305839
rect -62 -306815 -56 -305839
rect -102 -306827 -56 -306815
rect 56 -305839 102 -305827
rect 56 -306815 62 -305839
rect 96 -306815 102 -305839
rect 56 -306827 102 -306815
rect -46 -306865 46 -306859
rect -46 -306899 -34 -306865
rect 34 -306899 46 -306865
rect -46 -306905 46 -306899
rect -46 -306973 46 -306967
rect -46 -307007 -34 -306973
rect 34 -307007 46 -306973
rect -46 -307013 46 -307007
rect -102 -307057 -56 -307045
rect -102 -308033 -96 -307057
rect -62 -308033 -56 -307057
rect -102 -308045 -56 -308033
rect 56 -307057 102 -307045
rect 56 -308033 62 -307057
rect 96 -308033 102 -307057
rect 56 -308045 102 -308033
rect -46 -308083 46 -308077
rect -46 -308117 -34 -308083
rect 34 -308117 46 -308083
rect -46 -308123 46 -308117
rect -46 -308191 46 -308185
rect -46 -308225 -34 -308191
rect 34 -308225 46 -308191
rect -46 -308231 46 -308225
rect -102 -308275 -56 -308263
rect -102 -309251 -96 -308275
rect -62 -309251 -56 -308275
rect -102 -309263 -56 -309251
rect 56 -308275 102 -308263
rect 56 -309251 62 -308275
rect 96 -309251 102 -308275
rect 56 -309263 102 -309251
rect -46 -309301 46 -309295
rect -46 -309335 -34 -309301
rect 34 -309335 46 -309301
rect -46 -309341 46 -309335
rect -46 -309409 46 -309403
rect -46 -309443 -34 -309409
rect 34 -309443 46 -309409
rect -46 -309449 46 -309443
rect -102 -309493 -56 -309481
rect -102 -310469 -96 -309493
rect -62 -310469 -56 -309493
rect -102 -310481 -56 -310469
rect 56 -309493 102 -309481
rect 56 -310469 62 -309493
rect 96 -310469 102 -309493
rect 56 -310481 102 -310469
rect -46 -310519 46 -310513
rect -46 -310553 -34 -310519
rect 34 -310553 46 -310519
rect -46 -310559 46 -310553
rect -46 -310627 46 -310621
rect -46 -310661 -34 -310627
rect 34 -310661 46 -310627
rect -46 -310667 46 -310661
rect -102 -310711 -56 -310699
rect -102 -311687 -96 -310711
rect -62 -311687 -56 -310711
rect -102 -311699 -56 -311687
rect 56 -310711 102 -310699
rect 56 -311687 62 -310711
rect 96 -311687 102 -310711
rect 56 -311699 102 -311687
rect -46 -311737 46 -311731
rect -46 -311771 -34 -311737
rect 34 -311771 46 -311737
rect -46 -311777 46 -311771
rect -46 -311845 46 -311839
rect -46 -311879 -34 -311845
rect 34 -311879 46 -311845
rect -46 -311885 46 -311879
rect -102 -311929 -56 -311917
rect -102 -312905 -96 -311929
rect -62 -312905 -56 -311929
rect -102 -312917 -56 -312905
rect 56 -311929 102 -311917
rect 56 -312905 62 -311929
rect 96 -312905 102 -311929
rect 56 -312917 102 -312905
rect -46 -312955 46 -312949
rect -46 -312989 -34 -312955
rect 34 -312989 46 -312955
rect -46 -312995 46 -312989
rect -46 -313063 46 -313057
rect -46 -313097 -34 -313063
rect 34 -313097 46 -313063
rect -46 -313103 46 -313097
rect -102 -313147 -56 -313135
rect -102 -314123 -96 -313147
rect -62 -314123 -56 -313147
rect -102 -314135 -56 -314123
rect 56 -313147 102 -313135
rect 56 -314123 62 -313147
rect 96 -314123 102 -313147
rect 56 -314135 102 -314123
rect -46 -314173 46 -314167
rect -46 -314207 -34 -314173
rect 34 -314207 46 -314173
rect -46 -314213 46 -314207
rect -46 -314281 46 -314275
rect -46 -314315 -34 -314281
rect 34 -314315 46 -314281
rect -46 -314321 46 -314315
rect -102 -314365 -56 -314353
rect -102 -315341 -96 -314365
rect -62 -315341 -56 -314365
rect -102 -315353 -56 -315341
rect 56 -314365 102 -314353
rect 56 -315341 62 -314365
rect 96 -315341 102 -314365
rect 56 -315353 102 -315341
rect -46 -315391 46 -315385
rect -46 -315425 -34 -315391
rect 34 -315425 46 -315391
rect -46 -315431 46 -315425
rect -46 -315499 46 -315493
rect -46 -315533 -34 -315499
rect 34 -315533 46 -315499
rect -46 -315539 46 -315533
rect -102 -315583 -56 -315571
rect -102 -316559 -96 -315583
rect -62 -316559 -56 -315583
rect -102 -316571 -56 -316559
rect 56 -315583 102 -315571
rect 56 -316559 62 -315583
rect 96 -316559 102 -315583
rect 56 -316571 102 -316559
rect -46 -316609 46 -316603
rect -46 -316643 -34 -316609
rect 34 -316643 46 -316609
rect -46 -316649 46 -316643
rect -46 -316717 46 -316711
rect -46 -316751 -34 -316717
rect 34 -316751 46 -316717
rect -46 -316757 46 -316751
rect -102 -316801 -56 -316789
rect -102 -317777 -96 -316801
rect -62 -317777 -56 -316801
rect -102 -317789 -56 -317777
rect 56 -316801 102 -316789
rect 56 -317777 62 -316801
rect 96 -317777 102 -316801
rect 56 -317789 102 -317777
rect -46 -317827 46 -317821
rect -46 -317861 -34 -317827
rect 34 -317861 46 -317827
rect -46 -317867 46 -317861
rect -46 -317935 46 -317929
rect -46 -317969 -34 -317935
rect 34 -317969 46 -317935
rect -46 -317975 46 -317969
rect -102 -318019 -56 -318007
rect -102 -318995 -96 -318019
rect -62 -318995 -56 -318019
rect -102 -319007 -56 -318995
rect 56 -318019 102 -318007
rect 56 -318995 62 -318019
rect 96 -318995 102 -318019
rect 56 -319007 102 -318995
rect -46 -319045 46 -319039
rect -46 -319079 -34 -319045
rect 34 -319079 46 -319045
rect -46 -319085 46 -319079
rect -46 -319153 46 -319147
rect -46 -319187 -34 -319153
rect 34 -319187 46 -319153
rect -46 -319193 46 -319187
rect -102 -319237 -56 -319225
rect -102 -320213 -96 -319237
rect -62 -320213 -56 -319237
rect -102 -320225 -56 -320213
rect 56 -319237 102 -319225
rect 56 -320213 62 -319237
rect 96 -320213 102 -319237
rect 56 -320225 102 -320213
rect -46 -320263 46 -320257
rect -46 -320297 -34 -320263
rect 34 -320297 46 -320263
rect -46 -320303 46 -320297
rect -46 -320371 46 -320365
rect -46 -320405 -34 -320371
rect 34 -320405 46 -320371
rect -46 -320411 46 -320405
rect -102 -320455 -56 -320443
rect -102 -321431 -96 -320455
rect -62 -321431 -56 -320455
rect -102 -321443 -56 -321431
rect 56 -320455 102 -320443
rect 56 -321431 62 -320455
rect 96 -321431 102 -320455
rect 56 -321443 102 -321431
rect -46 -321481 46 -321475
rect -46 -321515 -34 -321481
rect 34 -321515 46 -321481
rect -46 -321521 46 -321515
rect -46 -321589 46 -321583
rect -46 -321623 -34 -321589
rect 34 -321623 46 -321589
rect -46 -321629 46 -321623
rect -102 -321673 -56 -321661
rect -102 -322649 -96 -321673
rect -62 -322649 -56 -321673
rect -102 -322661 -56 -322649
rect 56 -321673 102 -321661
rect 56 -322649 62 -321673
rect 96 -322649 102 -321673
rect 56 -322661 102 -322649
rect -46 -322699 46 -322693
rect -46 -322733 -34 -322699
rect 34 -322733 46 -322699
rect -46 -322739 46 -322733
rect -46 -322807 46 -322801
rect -46 -322841 -34 -322807
rect 34 -322841 46 -322807
rect -46 -322847 46 -322841
rect -102 -322891 -56 -322879
rect -102 -323867 -96 -322891
rect -62 -323867 -56 -322891
rect -102 -323879 -56 -323867
rect 56 -322891 102 -322879
rect 56 -323867 62 -322891
rect 96 -323867 102 -322891
rect 56 -323879 102 -323867
rect -46 -323917 46 -323911
rect -46 -323951 -34 -323917
rect 34 -323951 46 -323917
rect -46 -323957 46 -323951
rect -46 -324025 46 -324019
rect -46 -324059 -34 -324025
rect 34 -324059 46 -324025
rect -46 -324065 46 -324059
rect -102 -324109 -56 -324097
rect -102 -325085 -96 -324109
rect -62 -325085 -56 -324109
rect -102 -325097 -56 -325085
rect 56 -324109 102 -324097
rect 56 -325085 62 -324109
rect 96 -325085 102 -324109
rect 56 -325097 102 -325085
rect -46 -325135 46 -325129
rect -46 -325169 -34 -325135
rect 34 -325169 46 -325135
rect -46 -325175 46 -325169
rect -46 -325243 46 -325237
rect -46 -325277 -34 -325243
rect 34 -325277 46 -325243
rect -46 -325283 46 -325277
rect -102 -325327 -56 -325315
rect -102 -326303 -96 -325327
rect -62 -326303 -56 -325327
rect -102 -326315 -56 -326303
rect 56 -325327 102 -325315
rect 56 -326303 62 -325327
rect 96 -326303 102 -325327
rect 56 -326315 102 -326303
rect -46 -326353 46 -326347
rect -46 -326387 -34 -326353
rect 34 -326387 46 -326353
rect -46 -326393 46 -326387
rect -46 -326461 46 -326455
rect -46 -326495 -34 -326461
rect 34 -326495 46 -326461
rect -46 -326501 46 -326495
rect -102 -326545 -56 -326533
rect -102 -327521 -96 -326545
rect -62 -327521 -56 -326545
rect -102 -327533 -56 -327521
rect 56 -326545 102 -326533
rect 56 -327521 62 -326545
rect 96 -327521 102 -326545
rect 56 -327533 102 -327521
rect -46 -327571 46 -327565
rect -46 -327605 -34 -327571
rect 34 -327605 46 -327571
rect -46 -327611 46 -327605
rect -46 -327679 46 -327673
rect -46 -327713 -34 -327679
rect 34 -327713 46 -327679
rect -46 -327719 46 -327713
rect -102 -327763 -56 -327751
rect -102 -328739 -96 -327763
rect -62 -328739 -56 -327763
rect -102 -328751 -56 -328739
rect 56 -327763 102 -327751
rect 56 -328739 62 -327763
rect 96 -328739 102 -327763
rect 56 -328751 102 -328739
rect -46 -328789 46 -328783
rect -46 -328823 -34 -328789
rect 34 -328823 46 -328789
rect -46 -328829 46 -328823
rect -46 -328897 46 -328891
rect -46 -328931 -34 -328897
rect 34 -328931 46 -328897
rect -46 -328937 46 -328931
rect -102 -328981 -56 -328969
rect -102 -329957 -96 -328981
rect -62 -329957 -56 -328981
rect -102 -329969 -56 -329957
rect 56 -328981 102 -328969
rect 56 -329957 62 -328981
rect 96 -329957 102 -328981
rect 56 -329969 102 -329957
rect -46 -330007 46 -330001
rect -46 -330041 -34 -330007
rect 34 -330041 46 -330007
rect -46 -330047 46 -330041
rect -46 -330115 46 -330109
rect -46 -330149 -34 -330115
rect 34 -330149 46 -330115
rect -46 -330155 46 -330149
rect -102 -330199 -56 -330187
rect -102 -331175 -96 -330199
rect -62 -331175 -56 -330199
rect -102 -331187 -56 -331175
rect 56 -330199 102 -330187
rect 56 -331175 62 -330199
rect 96 -331175 102 -330199
rect 56 -331187 102 -331175
rect -46 -331225 46 -331219
rect -46 -331259 -34 -331225
rect 34 -331259 46 -331225
rect -46 -331265 46 -331259
rect -46 -331333 46 -331327
rect -46 -331367 -34 -331333
rect 34 -331367 46 -331333
rect -46 -331373 46 -331367
rect -102 -331417 -56 -331405
rect -102 -332393 -96 -331417
rect -62 -332393 -56 -331417
rect -102 -332405 -56 -332393
rect 56 -331417 102 -331405
rect 56 -332393 62 -331417
rect 96 -332393 102 -331417
rect 56 -332405 102 -332393
rect -46 -332443 46 -332437
rect -46 -332477 -34 -332443
rect 34 -332477 46 -332443
rect -46 -332483 46 -332477
rect -46 -332551 46 -332545
rect -46 -332585 -34 -332551
rect 34 -332585 46 -332551
rect -46 -332591 46 -332585
rect -102 -332635 -56 -332623
rect -102 -333611 -96 -332635
rect -62 -333611 -56 -332635
rect -102 -333623 -56 -333611
rect 56 -332635 102 -332623
rect 56 -333611 62 -332635
rect 96 -333611 102 -332635
rect 56 -333623 102 -333611
rect -46 -333661 46 -333655
rect -46 -333695 -34 -333661
rect 34 -333695 46 -333661
rect -46 -333701 46 -333695
rect -46 -333769 46 -333763
rect -46 -333803 -34 -333769
rect 34 -333803 46 -333769
rect -46 -333809 46 -333803
rect -102 -333853 -56 -333841
rect -102 -334829 -96 -333853
rect -62 -334829 -56 -333853
rect -102 -334841 -56 -334829
rect 56 -333853 102 -333841
rect 56 -334829 62 -333853
rect 96 -334829 102 -333853
rect 56 -334841 102 -334829
rect -46 -334879 46 -334873
rect -46 -334913 -34 -334879
rect 34 -334913 46 -334879
rect -46 -334919 46 -334913
rect -46 -334987 46 -334981
rect -46 -335021 -34 -334987
rect 34 -335021 46 -334987
rect -46 -335027 46 -335021
rect -102 -335071 -56 -335059
rect -102 -336047 -96 -335071
rect -62 -336047 -56 -335071
rect -102 -336059 -56 -336047
rect 56 -335071 102 -335059
rect 56 -336047 62 -335071
rect 96 -336047 102 -335071
rect 56 -336059 102 -336047
rect -46 -336097 46 -336091
rect -46 -336131 -34 -336097
rect 34 -336131 46 -336097
rect -46 -336137 46 -336131
rect -46 -336205 46 -336199
rect -46 -336239 -34 -336205
rect 34 -336239 46 -336205
rect -46 -336245 46 -336239
rect -102 -336289 -56 -336277
rect -102 -337265 -96 -336289
rect -62 -337265 -56 -336289
rect -102 -337277 -56 -337265
rect 56 -336289 102 -336277
rect 56 -337265 62 -336289
rect 96 -337265 102 -336289
rect 56 -337277 102 -337265
rect -46 -337315 46 -337309
rect -46 -337349 -34 -337315
rect 34 -337349 46 -337315
rect -46 -337355 46 -337349
rect -46 -337423 46 -337417
rect -46 -337457 -34 -337423
rect 34 -337457 46 -337423
rect -46 -337463 46 -337457
rect -102 -337507 -56 -337495
rect -102 -338483 -96 -337507
rect -62 -338483 -56 -337507
rect -102 -338495 -56 -338483
rect 56 -337507 102 -337495
rect 56 -338483 62 -337507
rect 96 -338483 102 -337507
rect 56 -338495 102 -338483
rect -46 -338533 46 -338527
rect -46 -338567 -34 -338533
rect 34 -338567 46 -338533
rect -46 -338573 46 -338567
rect -46 -338641 46 -338635
rect -46 -338675 -34 -338641
rect 34 -338675 46 -338641
rect -46 -338681 46 -338675
rect -102 -338725 -56 -338713
rect -102 -339701 -96 -338725
rect -62 -339701 -56 -338725
rect -102 -339713 -56 -339701
rect 56 -338725 102 -338713
rect 56 -339701 62 -338725
rect 96 -339701 102 -338725
rect 56 -339713 102 -339701
rect -46 -339751 46 -339745
rect -46 -339785 -34 -339751
rect 34 -339785 46 -339751
rect -46 -339791 46 -339785
rect -46 -339859 46 -339853
rect -46 -339893 -34 -339859
rect 34 -339893 46 -339859
rect -46 -339899 46 -339893
rect -102 -339943 -56 -339931
rect -102 -340919 -96 -339943
rect -62 -340919 -56 -339943
rect -102 -340931 -56 -340919
rect 56 -339943 102 -339931
rect 56 -340919 62 -339943
rect 96 -340919 102 -339943
rect 56 -340931 102 -340919
rect -46 -340969 46 -340963
rect -46 -341003 -34 -340969
rect 34 -341003 46 -340969
rect -46 -341009 46 -341003
rect -46 -341077 46 -341071
rect -46 -341111 -34 -341077
rect 34 -341111 46 -341077
rect -46 -341117 46 -341111
rect -102 -341161 -56 -341149
rect -102 -342137 -96 -341161
rect -62 -342137 -56 -341161
rect -102 -342149 -56 -342137
rect 56 -341161 102 -341149
rect 56 -342137 62 -341161
rect 96 -342137 102 -341161
rect 56 -342149 102 -342137
rect -46 -342187 46 -342181
rect -46 -342221 -34 -342187
rect 34 -342221 46 -342187
rect -46 -342227 46 -342221
rect -46 -342295 46 -342289
rect -46 -342329 -34 -342295
rect 34 -342329 46 -342295
rect -46 -342335 46 -342329
rect -102 -342379 -56 -342367
rect -102 -343355 -96 -342379
rect -62 -343355 -56 -342379
rect -102 -343367 -56 -343355
rect 56 -342379 102 -342367
rect 56 -343355 62 -342379
rect 96 -343355 102 -342379
rect 56 -343367 102 -343355
rect -46 -343405 46 -343399
rect -46 -343439 -34 -343405
rect 34 -343439 46 -343405
rect -46 -343445 46 -343439
rect -46 -343513 46 -343507
rect -46 -343547 -34 -343513
rect 34 -343547 46 -343513
rect -46 -343553 46 -343547
rect -102 -343597 -56 -343585
rect -102 -344573 -96 -343597
rect -62 -344573 -56 -343597
rect -102 -344585 -56 -344573
rect 56 -343597 102 -343585
rect 56 -344573 62 -343597
rect 96 -344573 102 -343597
rect 56 -344585 102 -344573
rect -46 -344623 46 -344617
rect -46 -344657 -34 -344623
rect 34 -344657 46 -344623
rect -46 -344663 46 -344657
rect -46 -344731 46 -344725
rect -46 -344765 -34 -344731
rect 34 -344765 46 -344731
rect -46 -344771 46 -344765
rect -102 -344815 -56 -344803
rect -102 -345791 -96 -344815
rect -62 -345791 -56 -344815
rect -102 -345803 -56 -345791
rect 56 -344815 102 -344803
rect 56 -345791 62 -344815
rect 96 -345791 102 -344815
rect 56 -345803 102 -345791
rect -46 -345841 46 -345835
rect -46 -345875 -34 -345841
rect 34 -345875 46 -345841
rect -46 -345881 46 -345875
rect -46 -345949 46 -345943
rect -46 -345983 -34 -345949
rect 34 -345983 46 -345949
rect -46 -345989 46 -345983
rect -102 -346033 -56 -346021
rect -102 -347009 -96 -346033
rect -62 -347009 -56 -346033
rect -102 -347021 -56 -347009
rect 56 -346033 102 -346021
rect 56 -347009 62 -346033
rect 96 -347009 102 -346033
rect 56 -347021 102 -347009
rect -46 -347059 46 -347053
rect -46 -347093 -34 -347059
rect 34 -347093 46 -347059
rect -46 -347099 46 -347093
rect -46 -347167 46 -347161
rect -46 -347201 -34 -347167
rect 34 -347201 46 -347167
rect -46 -347207 46 -347201
rect -102 -347251 -56 -347239
rect -102 -348227 -96 -347251
rect -62 -348227 -56 -347251
rect -102 -348239 -56 -348227
rect 56 -347251 102 -347239
rect 56 -348227 62 -347251
rect 96 -348227 102 -347251
rect 56 -348239 102 -348227
rect -46 -348277 46 -348271
rect -46 -348311 -34 -348277
rect 34 -348311 46 -348277
rect -46 -348317 46 -348311
rect -46 -348385 46 -348379
rect -46 -348419 -34 -348385
rect 34 -348419 46 -348385
rect -46 -348425 46 -348419
rect -102 -348469 -56 -348457
rect -102 -349445 -96 -348469
rect -62 -349445 -56 -348469
rect -102 -349457 -56 -349445
rect 56 -348469 102 -348457
rect 56 -349445 62 -348469
rect 96 -349445 102 -348469
rect 56 -349457 102 -349445
rect -46 -349495 46 -349489
rect -46 -349529 -34 -349495
rect 34 -349529 46 -349495
rect -46 -349535 46 -349529
rect -46 -349603 46 -349597
rect -46 -349637 -34 -349603
rect 34 -349637 46 -349603
rect -46 -349643 46 -349637
rect -102 -349687 -56 -349675
rect -102 -350663 -96 -349687
rect -62 -350663 -56 -349687
rect -102 -350675 -56 -350663
rect 56 -349687 102 -349675
rect 56 -350663 62 -349687
rect 96 -350663 102 -349687
rect 56 -350675 102 -350663
rect -46 -350713 46 -350707
rect -46 -350747 -34 -350713
rect 34 -350747 46 -350713
rect -46 -350753 46 -350747
rect -46 -350821 46 -350815
rect -46 -350855 -34 -350821
rect 34 -350855 46 -350821
rect -46 -350861 46 -350855
rect -102 -350905 -56 -350893
rect -102 -351881 -96 -350905
rect -62 -351881 -56 -350905
rect -102 -351893 -56 -351881
rect 56 -350905 102 -350893
rect 56 -351881 62 -350905
rect 96 -351881 102 -350905
rect 56 -351893 102 -351881
rect -46 -351931 46 -351925
rect -46 -351965 -34 -351931
rect 34 -351965 46 -351931
rect -46 -351971 46 -351965
rect -46 -352039 46 -352033
rect -46 -352073 -34 -352039
rect 34 -352073 46 -352039
rect -46 -352079 46 -352073
rect -102 -352123 -56 -352111
rect -102 -353099 -96 -352123
rect -62 -353099 -56 -352123
rect -102 -353111 -56 -353099
rect 56 -352123 102 -352111
rect 56 -353099 62 -352123
rect 96 -353099 102 -352123
rect 56 -353111 102 -353099
rect -46 -353149 46 -353143
rect -46 -353183 -34 -353149
rect 34 -353183 46 -353149
rect -46 -353189 46 -353183
rect -46 -353257 46 -353251
rect -46 -353291 -34 -353257
rect 34 -353291 46 -353257
rect -46 -353297 46 -353291
rect -102 -353341 -56 -353329
rect -102 -354317 -96 -353341
rect -62 -354317 -56 -353341
rect -102 -354329 -56 -354317
rect 56 -353341 102 -353329
rect 56 -354317 62 -353341
rect 96 -354317 102 -353341
rect 56 -354329 102 -354317
rect -46 -354367 46 -354361
rect -46 -354401 -34 -354367
rect 34 -354401 46 -354367
rect -46 -354407 46 -354401
rect -46 -354475 46 -354469
rect -46 -354509 -34 -354475
rect 34 -354509 46 -354475
rect -46 -354515 46 -354509
rect -102 -354559 -56 -354547
rect -102 -355535 -96 -354559
rect -62 -355535 -56 -354559
rect -102 -355547 -56 -355535
rect 56 -354559 102 -354547
rect 56 -355535 62 -354559
rect 96 -355535 102 -354559
rect 56 -355547 102 -355535
rect -46 -355585 46 -355579
rect -46 -355619 -34 -355585
rect 34 -355619 46 -355585
rect -46 -355625 46 -355619
rect -46 -355693 46 -355687
rect -46 -355727 -34 -355693
rect 34 -355727 46 -355693
rect -46 -355733 46 -355727
rect -102 -355777 -56 -355765
rect -102 -356753 -96 -355777
rect -62 -356753 -56 -355777
rect -102 -356765 -56 -356753
rect 56 -355777 102 -355765
rect 56 -356753 62 -355777
rect 96 -356753 102 -355777
rect 56 -356765 102 -356753
rect -46 -356803 46 -356797
rect -46 -356837 -34 -356803
rect 34 -356837 46 -356803
rect -46 -356843 46 -356837
rect -46 -356911 46 -356905
rect -46 -356945 -34 -356911
rect 34 -356945 46 -356911
rect -46 -356951 46 -356945
rect -102 -356995 -56 -356983
rect -102 -357971 -96 -356995
rect -62 -357971 -56 -356995
rect -102 -357983 -56 -357971
rect 56 -356995 102 -356983
rect 56 -357971 62 -356995
rect 96 -357971 102 -356995
rect 56 -357983 102 -357971
rect -46 -358021 46 -358015
rect -46 -358055 -34 -358021
rect 34 -358055 46 -358021
rect -46 -358061 46 -358055
rect -46 -358129 46 -358123
rect -46 -358163 -34 -358129
rect 34 -358163 46 -358129
rect -46 -358169 46 -358163
rect -102 -358213 -56 -358201
rect -102 -359189 -96 -358213
rect -62 -359189 -56 -358213
rect -102 -359201 -56 -359189
rect 56 -358213 102 -358201
rect 56 -359189 62 -358213
rect 96 -359189 102 -358213
rect 56 -359201 102 -359189
rect -46 -359239 46 -359233
rect -46 -359273 -34 -359239
rect 34 -359273 46 -359239
rect -46 -359279 46 -359273
rect -46 -359347 46 -359341
rect -46 -359381 -34 -359347
rect 34 -359381 46 -359347
rect -46 -359387 46 -359381
rect -102 -359431 -56 -359419
rect -102 -360407 -96 -359431
rect -62 -360407 -56 -359431
rect -102 -360419 -56 -360407
rect 56 -359431 102 -359419
rect 56 -360407 62 -359431
rect 96 -360407 102 -359431
rect 56 -360419 102 -360407
rect -46 -360457 46 -360451
rect -46 -360491 -34 -360457
rect 34 -360491 46 -360457
rect -46 -360497 46 -360491
rect -46 -360565 46 -360559
rect -46 -360599 -34 -360565
rect 34 -360599 46 -360565
rect -46 -360605 46 -360599
rect -102 -360649 -56 -360637
rect -102 -361625 -96 -360649
rect -62 -361625 -56 -360649
rect -102 -361637 -56 -361625
rect 56 -360649 102 -360637
rect 56 -361625 62 -360649
rect 96 -361625 102 -360649
rect 56 -361637 102 -361625
rect -46 -361675 46 -361669
rect -46 -361709 -34 -361675
rect 34 -361709 46 -361675
rect -46 -361715 46 -361709
rect -46 -361783 46 -361777
rect -46 -361817 -34 -361783
rect 34 -361817 46 -361783
rect -46 -361823 46 -361817
rect -102 -361867 -56 -361855
rect -102 -362843 -96 -361867
rect -62 -362843 -56 -361867
rect -102 -362855 -56 -362843
rect 56 -361867 102 -361855
rect 56 -362843 62 -361867
rect 96 -362843 102 -361867
rect 56 -362855 102 -362843
rect -46 -362893 46 -362887
rect -46 -362927 -34 -362893
rect 34 -362927 46 -362893
rect -46 -362933 46 -362927
rect -46 -363001 46 -362995
rect -46 -363035 -34 -363001
rect 34 -363035 46 -363001
rect -46 -363041 46 -363035
rect -102 -363085 -56 -363073
rect -102 -364061 -96 -363085
rect -62 -364061 -56 -363085
rect -102 -364073 -56 -364061
rect 56 -363085 102 -363073
rect 56 -364061 62 -363085
rect 96 -364061 102 -363085
rect 56 -364073 102 -364061
rect -46 -364111 46 -364105
rect -46 -364145 -34 -364111
rect 34 -364145 46 -364111
rect -46 -364151 46 -364145
rect -46 -364219 46 -364213
rect -46 -364253 -34 -364219
rect 34 -364253 46 -364219
rect -46 -364259 46 -364253
rect -102 -364303 -56 -364291
rect -102 -365279 -96 -364303
rect -62 -365279 -56 -364303
rect -102 -365291 -56 -365279
rect 56 -364303 102 -364291
rect 56 -365279 62 -364303
rect 96 -365279 102 -364303
rect 56 -365291 102 -365279
rect -46 -365329 46 -365323
rect -46 -365363 -34 -365329
rect 34 -365363 46 -365329
rect -46 -365369 46 -365363
rect -46 -365437 46 -365431
rect -46 -365471 -34 -365437
rect 34 -365471 46 -365437
rect -46 -365477 46 -365471
rect -102 -365521 -56 -365509
rect -102 -366497 -96 -365521
rect -62 -366497 -56 -365521
rect -102 -366509 -56 -366497
rect 56 -365521 102 -365509
rect 56 -366497 62 -365521
rect 96 -366497 102 -365521
rect 56 -366509 102 -366497
rect -46 -366547 46 -366541
rect -46 -366581 -34 -366547
rect 34 -366581 46 -366547
rect -46 -366587 46 -366581
rect -46 -366655 46 -366649
rect -46 -366689 -34 -366655
rect 34 -366689 46 -366655
rect -46 -366695 46 -366689
rect -102 -366739 -56 -366727
rect -102 -367715 -96 -366739
rect -62 -367715 -56 -366739
rect -102 -367727 -56 -367715
rect 56 -366739 102 -366727
rect 56 -367715 62 -366739
rect 96 -367715 102 -366739
rect 56 -367727 102 -367715
rect -46 -367765 46 -367759
rect -46 -367799 -34 -367765
rect 34 -367799 46 -367765
rect -46 -367805 46 -367799
rect -46 -367873 46 -367867
rect -46 -367907 -34 -367873
rect 34 -367907 46 -367873
rect -46 -367913 46 -367907
rect -102 -367957 -56 -367945
rect -102 -368933 -96 -367957
rect -62 -368933 -56 -367957
rect -102 -368945 -56 -368933
rect 56 -367957 102 -367945
rect 56 -368933 62 -367957
rect 96 -368933 102 -367957
rect 56 -368945 102 -368933
rect -46 -368983 46 -368977
rect -46 -369017 -34 -368983
rect 34 -369017 46 -368983
rect -46 -369023 46 -369017
rect -46 -369091 46 -369085
rect -46 -369125 -34 -369091
rect 34 -369125 46 -369091
rect -46 -369131 46 -369125
rect -102 -369175 -56 -369163
rect -102 -370151 -96 -369175
rect -62 -370151 -56 -369175
rect -102 -370163 -56 -370151
rect 56 -369175 102 -369163
rect 56 -370151 62 -369175
rect 96 -370151 102 -369175
rect 56 -370163 102 -370151
rect -46 -370201 46 -370195
rect -46 -370235 -34 -370201
rect 34 -370235 46 -370201
rect -46 -370241 46 -370235
rect -46 -370309 46 -370303
rect -46 -370343 -34 -370309
rect 34 -370343 46 -370309
rect -46 -370349 46 -370343
rect -102 -370393 -56 -370381
rect -102 -371369 -96 -370393
rect -62 -371369 -56 -370393
rect -102 -371381 -56 -371369
rect 56 -370393 102 -370381
rect 56 -371369 62 -370393
rect 96 -371369 102 -370393
rect 56 -371381 102 -371369
rect -46 -371419 46 -371413
rect -46 -371453 -34 -371419
rect 34 -371453 46 -371419
rect -46 -371459 46 -371453
rect -46 -371527 46 -371521
rect -46 -371561 -34 -371527
rect 34 -371561 46 -371527
rect -46 -371567 46 -371561
rect -102 -371611 -56 -371599
rect -102 -372587 -96 -371611
rect -62 -372587 -56 -371611
rect -102 -372599 -56 -372587
rect 56 -371611 102 -371599
rect 56 -372587 62 -371611
rect 96 -372587 102 -371611
rect 56 -372599 102 -372587
rect -46 -372637 46 -372631
rect -46 -372671 -34 -372637
rect 34 -372671 46 -372637
rect -46 -372677 46 -372671
rect -46 -372745 46 -372739
rect -46 -372779 -34 -372745
rect 34 -372779 46 -372745
rect -46 -372785 46 -372779
rect -102 -372829 -56 -372817
rect -102 -373805 -96 -372829
rect -62 -373805 -56 -372829
rect -102 -373817 -56 -373805
rect 56 -372829 102 -372817
rect 56 -373805 62 -372829
rect 96 -373805 102 -372829
rect 56 -373817 102 -373805
rect -46 -373855 46 -373849
rect -46 -373889 -34 -373855
rect 34 -373889 46 -373855
rect -46 -373895 46 -373889
rect -46 -373963 46 -373957
rect -46 -373997 -34 -373963
rect 34 -373997 46 -373963
rect -46 -374003 46 -373997
rect -102 -374047 -56 -374035
rect -102 -375023 -96 -374047
rect -62 -375023 -56 -374047
rect -102 -375035 -56 -375023
rect 56 -374047 102 -374035
rect 56 -375023 62 -374047
rect 96 -375023 102 -374047
rect 56 -375035 102 -375023
rect -46 -375073 46 -375067
rect -46 -375107 -34 -375073
rect 34 -375107 46 -375073
rect -46 -375113 46 -375107
rect -46 -375181 46 -375175
rect -46 -375215 -34 -375181
rect 34 -375215 46 -375181
rect -46 -375221 46 -375215
rect -102 -375265 -56 -375253
rect -102 -376241 -96 -375265
rect -62 -376241 -56 -375265
rect -102 -376253 -56 -376241
rect 56 -375265 102 -375253
rect 56 -376241 62 -375265
rect 96 -376241 102 -375265
rect 56 -376253 102 -376241
rect -46 -376291 46 -376285
rect -46 -376325 -34 -376291
rect 34 -376325 46 -376291
rect -46 -376331 46 -376325
rect -46 -376399 46 -376393
rect -46 -376433 -34 -376399
rect 34 -376433 46 -376399
rect -46 -376439 46 -376433
rect -102 -376483 -56 -376471
rect -102 -377459 -96 -376483
rect -62 -377459 -56 -376483
rect -102 -377471 -56 -377459
rect 56 -376483 102 -376471
rect 56 -377459 62 -376483
rect 96 -377459 102 -376483
rect 56 -377471 102 -377459
rect -46 -377509 46 -377503
rect -46 -377543 -34 -377509
rect 34 -377543 46 -377509
rect -46 -377549 46 -377543
rect -46 -377617 46 -377611
rect -46 -377651 -34 -377617
rect 34 -377651 46 -377617
rect -46 -377657 46 -377651
rect -102 -377701 -56 -377689
rect -102 -378677 -96 -377701
rect -62 -378677 -56 -377701
rect -102 -378689 -56 -378677
rect 56 -377701 102 -377689
rect 56 -378677 62 -377701
rect 96 -378677 102 -377701
rect 56 -378689 102 -378677
rect -46 -378727 46 -378721
rect -46 -378761 -34 -378727
rect 34 -378761 46 -378727
rect -46 -378767 46 -378761
rect -46 -378835 46 -378829
rect -46 -378869 -34 -378835
rect 34 -378869 46 -378835
rect -46 -378875 46 -378869
rect -102 -378919 -56 -378907
rect -102 -379895 -96 -378919
rect -62 -379895 -56 -378919
rect -102 -379907 -56 -379895
rect 56 -378919 102 -378907
rect 56 -379895 62 -378919
rect 96 -379895 102 -378919
rect 56 -379907 102 -379895
rect -46 -379945 46 -379939
rect -46 -379979 -34 -379945
rect 34 -379979 46 -379945
rect -46 -379985 46 -379979
rect -46 -380053 46 -380047
rect -46 -380087 -34 -380053
rect 34 -380087 46 -380053
rect -46 -380093 46 -380087
rect -102 -380137 -56 -380125
rect -102 -381113 -96 -380137
rect -62 -381113 -56 -380137
rect -102 -381125 -56 -381113
rect 56 -380137 102 -380125
rect 56 -381113 62 -380137
rect 96 -381113 102 -380137
rect 56 -381125 102 -381113
rect -46 -381163 46 -381157
rect -46 -381197 -34 -381163
rect 34 -381197 46 -381163
rect -46 -381203 46 -381197
rect -46 -381271 46 -381265
rect -46 -381305 -34 -381271
rect 34 -381305 46 -381271
rect -46 -381311 46 -381305
rect -102 -381355 -56 -381343
rect -102 -382331 -96 -381355
rect -62 -382331 -56 -381355
rect -102 -382343 -56 -382331
rect 56 -381355 102 -381343
rect 56 -382331 62 -381355
rect 96 -382331 102 -381355
rect 56 -382343 102 -382331
rect -46 -382381 46 -382375
rect -46 -382415 -34 -382381
rect 34 -382415 46 -382381
rect -46 -382421 46 -382415
rect -46 -382489 46 -382483
rect -46 -382523 -34 -382489
rect 34 -382523 46 -382489
rect -46 -382529 46 -382523
rect -102 -382573 -56 -382561
rect -102 -383549 -96 -382573
rect -62 -383549 -56 -382573
rect -102 -383561 -56 -383549
rect 56 -382573 102 -382561
rect 56 -383549 62 -382573
rect 96 -383549 102 -382573
rect 56 -383561 102 -383549
rect -46 -383599 46 -383593
rect -46 -383633 -34 -383599
rect 34 -383633 46 -383599
rect -46 -383639 46 -383633
rect -46 -383707 46 -383701
rect -46 -383741 -34 -383707
rect 34 -383741 46 -383707
rect -46 -383747 46 -383741
rect -102 -383791 -56 -383779
rect -102 -384767 -96 -383791
rect -62 -384767 -56 -383791
rect -102 -384779 -56 -384767
rect 56 -383791 102 -383779
rect 56 -384767 62 -383791
rect 96 -384767 102 -383791
rect 56 -384779 102 -384767
rect -46 -384817 46 -384811
rect -46 -384851 -34 -384817
rect 34 -384851 46 -384817
rect -46 -384857 46 -384851
rect -46 -384925 46 -384919
rect -46 -384959 -34 -384925
rect 34 -384959 46 -384925
rect -46 -384965 46 -384959
rect -102 -385009 -56 -384997
rect -102 -385985 -96 -385009
rect -62 -385985 -56 -385009
rect -102 -385997 -56 -385985
rect 56 -385009 102 -384997
rect 56 -385985 62 -385009
rect 96 -385985 102 -385009
rect 56 -385997 102 -385985
rect -46 -386035 46 -386029
rect -46 -386069 -34 -386035
rect 34 -386069 46 -386035
rect -46 -386075 46 -386069
rect -46 -386143 46 -386137
rect -46 -386177 -34 -386143
rect 34 -386177 46 -386143
rect -46 -386183 46 -386177
rect -102 -386227 -56 -386215
rect -102 -387203 -96 -386227
rect -62 -387203 -56 -386227
rect -102 -387215 -56 -387203
rect 56 -386227 102 -386215
rect 56 -387203 62 -386227
rect 96 -387203 102 -386227
rect 56 -387215 102 -387203
rect -46 -387253 46 -387247
rect -46 -387287 -34 -387253
rect 34 -387287 46 -387253
rect -46 -387293 46 -387287
rect -46 -387361 46 -387355
rect -46 -387395 -34 -387361
rect 34 -387395 46 -387361
rect -46 -387401 46 -387395
rect -102 -387445 -56 -387433
rect -102 -388421 -96 -387445
rect -62 -388421 -56 -387445
rect -102 -388433 -56 -388421
rect 56 -387445 102 -387433
rect 56 -388421 62 -387445
rect 96 -388421 102 -387445
rect 56 -388433 102 -388421
rect -46 -388471 46 -388465
rect -46 -388505 -34 -388471
rect 34 -388505 46 -388471
rect -46 -388511 46 -388505
rect -46 -388579 46 -388573
rect -46 -388613 -34 -388579
rect 34 -388613 46 -388579
rect -46 -388619 46 -388613
rect -102 -388663 -56 -388651
rect -102 -389639 -96 -388663
rect -62 -389639 -56 -388663
rect -102 -389651 -56 -389639
rect 56 -388663 102 -388651
rect 56 -389639 62 -388663
rect 96 -389639 102 -388663
rect 56 -389651 102 -389639
rect -46 -389689 46 -389683
rect -46 -389723 -34 -389689
rect 34 -389723 46 -389689
rect -46 -389729 46 -389723
rect -46 -389797 46 -389791
rect -46 -389831 -34 -389797
rect 34 -389831 46 -389797
rect -46 -389837 46 -389831
rect -102 -389881 -56 -389869
rect -102 -390857 -96 -389881
rect -62 -390857 -56 -389881
rect -102 -390869 -56 -390857
rect 56 -389881 102 -389869
rect 56 -390857 62 -389881
rect 96 -390857 102 -389881
rect 56 -390869 102 -390857
rect -46 -390907 46 -390901
rect -46 -390941 -34 -390907
rect 34 -390941 46 -390907
rect -46 -390947 46 -390941
rect -46 -391015 46 -391009
rect -46 -391049 -34 -391015
rect 34 -391049 46 -391015
rect -46 -391055 46 -391049
rect -102 -391099 -56 -391087
rect -102 -392075 -96 -391099
rect -62 -392075 -56 -391099
rect -102 -392087 -56 -392075
rect 56 -391099 102 -391087
rect 56 -392075 62 -391099
rect 96 -392075 102 -391099
rect 56 -392087 102 -392075
rect -46 -392125 46 -392119
rect -46 -392159 -34 -392125
rect 34 -392159 46 -392125
rect -46 -392165 46 -392159
rect -46 -392233 46 -392227
rect -46 -392267 -34 -392233
rect 34 -392267 46 -392233
rect -46 -392273 46 -392267
rect -102 -392317 -56 -392305
rect -102 -393293 -96 -392317
rect -62 -393293 -56 -392317
rect -102 -393305 -56 -393293
rect 56 -392317 102 -392305
rect 56 -393293 62 -392317
rect 96 -393293 102 -392317
rect 56 -393305 102 -393293
rect -46 -393343 46 -393337
rect -46 -393377 -34 -393343
rect 34 -393377 46 -393343
rect -46 -393383 46 -393377
rect -46 -393451 46 -393445
rect -46 -393485 -34 -393451
rect 34 -393485 46 -393451
rect -46 -393491 46 -393485
rect -102 -393535 -56 -393523
rect -102 -394511 -96 -393535
rect -62 -394511 -56 -393535
rect -102 -394523 -56 -394511
rect 56 -393535 102 -393523
rect 56 -394511 62 -393535
rect 96 -394511 102 -393535
rect 56 -394523 102 -394511
rect -46 -394561 46 -394555
rect -46 -394595 -34 -394561
rect 34 -394595 46 -394561
rect -46 -394601 46 -394595
rect -46 -394669 46 -394663
rect -46 -394703 -34 -394669
rect 34 -394703 46 -394669
rect -46 -394709 46 -394703
rect -102 -394753 -56 -394741
rect -102 -395729 -96 -394753
rect -62 -395729 -56 -394753
rect -102 -395741 -56 -395729
rect 56 -394753 102 -394741
rect 56 -395729 62 -394753
rect 96 -395729 102 -394753
rect 56 -395741 102 -395729
rect -46 -395779 46 -395773
rect -46 -395813 -34 -395779
rect 34 -395813 46 -395779
rect -46 -395819 46 -395813
rect -46 -395887 46 -395881
rect -46 -395921 -34 -395887
rect 34 -395921 46 -395887
rect -46 -395927 46 -395921
rect -102 -395971 -56 -395959
rect -102 -396947 -96 -395971
rect -62 -396947 -56 -395971
rect -102 -396959 -56 -396947
rect 56 -395971 102 -395959
rect 56 -396947 62 -395971
rect 96 -396947 102 -395971
rect 56 -396959 102 -396947
rect -46 -396997 46 -396991
rect -46 -397031 -34 -396997
rect 34 -397031 46 -396997
rect -46 -397037 46 -397031
rect -46 -397105 46 -397099
rect -46 -397139 -34 -397105
rect 34 -397139 46 -397105
rect -46 -397145 46 -397139
rect -102 -397189 -56 -397177
rect -102 -398165 -96 -397189
rect -62 -398165 -56 -397189
rect -102 -398177 -56 -398165
rect 56 -397189 102 -397177
rect 56 -398165 62 -397189
rect 96 -398165 102 -397189
rect 56 -398177 102 -398165
rect -46 -398215 46 -398209
rect -46 -398249 -34 -398215
rect 34 -398249 46 -398215
rect -46 -398255 46 -398249
rect -46 -398323 46 -398317
rect -46 -398357 -34 -398323
rect 34 -398357 46 -398323
rect -46 -398363 46 -398357
rect -102 -398407 -56 -398395
rect -102 -399383 -96 -398407
rect -62 -399383 -56 -398407
rect -102 -399395 -56 -399383
rect 56 -398407 102 -398395
rect 56 -399383 62 -398407
rect 96 -399383 102 -398407
rect 56 -399395 102 -399383
rect -46 -399433 46 -399427
rect -46 -399467 -34 -399433
rect 34 -399467 46 -399433
rect -46 -399473 46 -399467
rect -46 -399541 46 -399535
rect -46 -399575 -34 -399541
rect 34 -399575 46 -399541
rect -46 -399581 46 -399575
rect -102 -399625 -56 -399613
rect -102 -400601 -96 -399625
rect -62 -400601 -56 -399625
rect -102 -400613 -56 -400601
rect 56 -399625 102 -399613
rect 56 -400601 62 -399625
rect 96 -400601 102 -399625
rect 56 -400613 102 -400601
rect -46 -400651 46 -400645
rect -46 -400685 -34 -400651
rect 34 -400685 46 -400651
rect -46 -400691 46 -400685
rect -46 -400759 46 -400753
rect -46 -400793 -34 -400759
rect 34 -400793 46 -400759
rect -46 -400799 46 -400793
rect -102 -400843 -56 -400831
rect -102 -401819 -96 -400843
rect -62 -401819 -56 -400843
rect -102 -401831 -56 -401819
rect 56 -400843 102 -400831
rect 56 -401819 62 -400843
rect 96 -401819 102 -400843
rect 56 -401831 102 -401819
rect -46 -401869 46 -401863
rect -46 -401903 -34 -401869
rect 34 -401903 46 -401869
rect -46 -401909 46 -401903
rect -46 -401977 46 -401971
rect -46 -402011 -34 -401977
rect 34 -402011 46 -401977
rect -46 -402017 46 -402011
rect -102 -402061 -56 -402049
rect -102 -403037 -96 -402061
rect -62 -403037 -56 -402061
rect -102 -403049 -56 -403037
rect 56 -402061 102 -402049
rect 56 -403037 62 -402061
rect 96 -403037 102 -402061
rect 56 -403049 102 -403037
rect -46 -403087 46 -403081
rect -46 -403121 -34 -403087
rect 34 -403121 46 -403087
rect -46 -403127 46 -403121
rect -46 -403195 46 -403189
rect -46 -403229 -34 -403195
rect 34 -403229 46 -403195
rect -46 -403235 46 -403229
rect -102 -403279 -56 -403267
rect -102 -404255 -96 -403279
rect -62 -404255 -56 -403279
rect -102 -404267 -56 -404255
rect 56 -403279 102 -403267
rect 56 -404255 62 -403279
rect 96 -404255 102 -403279
rect 56 -404267 102 -404255
rect -46 -404305 46 -404299
rect -46 -404339 -34 -404305
rect 34 -404339 46 -404305
rect -46 -404345 46 -404339
rect -46 -404413 46 -404407
rect -46 -404447 -34 -404413
rect 34 -404447 46 -404413
rect -46 -404453 46 -404447
rect -102 -404497 -56 -404485
rect -102 -405473 -96 -404497
rect -62 -405473 -56 -404497
rect -102 -405485 -56 -405473
rect 56 -404497 102 -404485
rect 56 -405473 62 -404497
rect 96 -405473 102 -404497
rect 56 -405485 102 -405473
rect -46 -405523 46 -405517
rect -46 -405557 -34 -405523
rect 34 -405557 46 -405523
rect -46 -405563 46 -405557
rect -46 -405631 46 -405625
rect -46 -405665 -34 -405631
rect 34 -405665 46 -405631
rect -46 -405671 46 -405665
rect -102 -405715 -56 -405703
rect -102 -406691 -96 -405715
rect -62 -406691 -56 -405715
rect -102 -406703 -56 -406691
rect 56 -405715 102 -405703
rect 56 -406691 62 -405715
rect 96 -406691 102 -405715
rect 56 -406703 102 -406691
rect -46 -406741 46 -406735
rect -46 -406775 -34 -406741
rect 34 -406775 46 -406741
rect -46 -406781 46 -406775
rect -46 -406849 46 -406843
rect -46 -406883 -34 -406849
rect 34 -406883 46 -406849
rect -46 -406889 46 -406883
rect -102 -406933 -56 -406921
rect -102 -407909 -96 -406933
rect -62 -407909 -56 -406933
rect -102 -407921 -56 -407909
rect 56 -406933 102 -406921
rect 56 -407909 62 -406933
rect 96 -407909 102 -406933
rect 56 -407921 102 -407909
rect -46 -407959 46 -407953
rect -46 -407993 -34 -407959
rect 34 -407993 46 -407959
rect -46 -407999 46 -407993
rect -46 -408067 46 -408061
rect -46 -408101 -34 -408067
rect 34 -408101 46 -408067
rect -46 -408107 46 -408101
rect -102 -408151 -56 -408139
rect -102 -409127 -96 -408151
rect -62 -409127 -56 -408151
rect -102 -409139 -56 -409127
rect 56 -408151 102 -408139
rect 56 -409127 62 -408151
rect 96 -409127 102 -408151
rect 56 -409139 102 -409127
rect -46 -409177 46 -409171
rect -46 -409211 -34 -409177
rect 34 -409211 46 -409177
rect -46 -409217 46 -409211
rect -46 -409285 46 -409279
rect -46 -409319 -34 -409285
rect 34 -409319 46 -409285
rect -46 -409325 46 -409319
rect -102 -409369 -56 -409357
rect -102 -410345 -96 -409369
rect -62 -410345 -56 -409369
rect -102 -410357 -56 -410345
rect 56 -409369 102 -409357
rect 56 -410345 62 -409369
rect 96 -410345 102 -409369
rect 56 -410357 102 -410345
rect -46 -410395 46 -410389
rect -46 -410429 -34 -410395
rect 34 -410429 46 -410395
rect -46 -410435 46 -410429
rect -46 -410503 46 -410497
rect -46 -410537 -34 -410503
rect 34 -410537 46 -410503
rect -46 -410543 46 -410537
rect -102 -410587 -56 -410575
rect -102 -411563 -96 -410587
rect -62 -411563 -56 -410587
rect -102 -411575 -56 -411563
rect 56 -410587 102 -410575
rect 56 -411563 62 -410587
rect 96 -411563 102 -410587
rect 56 -411575 102 -411563
rect -46 -411613 46 -411607
rect -46 -411647 -34 -411613
rect 34 -411647 46 -411613
rect -46 -411653 46 -411647
rect -46 -411721 46 -411715
rect -46 -411755 -34 -411721
rect 34 -411755 46 -411721
rect -46 -411761 46 -411755
rect -102 -411805 -56 -411793
rect -102 -412781 -96 -411805
rect -62 -412781 -56 -411805
rect -102 -412793 -56 -412781
rect 56 -411805 102 -411793
rect 56 -412781 62 -411805
rect 96 -412781 102 -411805
rect 56 -412793 102 -412781
rect -46 -412831 46 -412825
rect -46 -412865 -34 -412831
rect 34 -412865 46 -412831
rect -46 -412871 46 -412865
rect -46 -412939 46 -412933
rect -46 -412973 -34 -412939
rect 34 -412973 46 -412939
rect -46 -412979 46 -412973
rect -102 -413023 -56 -413011
rect -102 -413999 -96 -413023
rect -62 -413999 -56 -413023
rect -102 -414011 -56 -413999
rect 56 -413023 102 -413011
rect 56 -413999 62 -413023
rect 96 -413999 102 -413023
rect 56 -414011 102 -413999
rect -46 -414049 46 -414043
rect -46 -414083 -34 -414049
rect 34 -414083 46 -414049
rect -46 -414089 46 -414083
rect -46 -414157 46 -414151
rect -46 -414191 -34 -414157
rect 34 -414191 46 -414157
rect -46 -414197 46 -414191
rect -102 -414241 -56 -414229
rect -102 -415217 -96 -414241
rect -62 -415217 -56 -414241
rect -102 -415229 -56 -415217
rect 56 -414241 102 -414229
rect 56 -415217 62 -414241
rect 96 -415217 102 -414241
rect 56 -415229 102 -415217
rect -46 -415267 46 -415261
rect -46 -415301 -34 -415267
rect 34 -415301 46 -415267
rect -46 -415307 46 -415301
rect -46 -415375 46 -415369
rect -46 -415409 -34 -415375
rect 34 -415409 46 -415375
rect -46 -415415 46 -415409
rect -102 -415459 -56 -415447
rect -102 -416435 -96 -415459
rect -62 -416435 -56 -415459
rect -102 -416447 -56 -416435
rect 56 -415459 102 -415447
rect 56 -416435 62 -415459
rect 96 -416435 102 -415459
rect 56 -416447 102 -416435
rect -46 -416485 46 -416479
rect -46 -416519 -34 -416485
rect 34 -416519 46 -416485
rect -46 -416525 46 -416519
rect -46 -416593 46 -416587
rect -46 -416627 -34 -416593
rect 34 -416627 46 -416593
rect -46 -416633 46 -416627
rect -102 -416677 -56 -416665
rect -102 -417653 -96 -416677
rect -62 -417653 -56 -416677
rect -102 -417665 -56 -417653
rect 56 -416677 102 -416665
rect 56 -417653 62 -416677
rect 96 -417653 102 -416677
rect 56 -417665 102 -417653
rect -46 -417703 46 -417697
rect -46 -417737 -34 -417703
rect 34 -417737 46 -417703
rect -46 -417743 46 -417737
rect -46 -417811 46 -417805
rect -46 -417845 -34 -417811
rect 34 -417845 46 -417811
rect -46 -417851 46 -417845
rect -102 -417895 -56 -417883
rect -102 -418871 -96 -417895
rect -62 -418871 -56 -417895
rect -102 -418883 -56 -418871
rect 56 -417895 102 -417883
rect 56 -418871 62 -417895
rect 96 -418871 102 -417895
rect 56 -418883 102 -418871
rect -46 -418921 46 -418915
rect -46 -418955 -34 -418921
rect 34 -418955 46 -418921
rect -46 -418961 46 -418955
rect -46 -419029 46 -419023
rect -46 -419063 -34 -419029
rect 34 -419063 46 -419029
rect -46 -419069 46 -419063
rect -102 -419113 -56 -419101
rect -102 -420089 -96 -419113
rect -62 -420089 -56 -419113
rect -102 -420101 -56 -420089
rect 56 -419113 102 -419101
rect 56 -420089 62 -419113
rect 96 -420089 102 -419113
rect 56 -420101 102 -420089
rect -46 -420139 46 -420133
rect -46 -420173 -34 -420139
rect 34 -420173 46 -420139
rect -46 -420179 46 -420173
rect -46 -420247 46 -420241
rect -46 -420281 -34 -420247
rect 34 -420281 46 -420247
rect -46 -420287 46 -420281
rect -102 -420331 -56 -420319
rect -102 -421307 -96 -420331
rect -62 -421307 -56 -420331
rect -102 -421319 -56 -421307
rect 56 -420331 102 -420319
rect 56 -421307 62 -420331
rect 96 -421307 102 -420331
rect 56 -421319 102 -421307
rect -46 -421357 46 -421351
rect -46 -421391 -34 -421357
rect 34 -421391 46 -421357
rect -46 -421397 46 -421391
rect -46 -421465 46 -421459
rect -46 -421499 -34 -421465
rect 34 -421499 46 -421465
rect -46 -421505 46 -421499
rect -102 -421549 -56 -421537
rect -102 -422525 -96 -421549
rect -62 -422525 -56 -421549
rect -102 -422537 -56 -422525
rect 56 -421549 102 -421537
rect 56 -422525 62 -421549
rect 96 -422525 102 -421549
rect 56 -422537 102 -422525
rect -46 -422575 46 -422569
rect -46 -422609 -34 -422575
rect 34 -422609 46 -422575
rect -46 -422615 46 -422609
rect -46 -422683 46 -422677
rect -46 -422717 -34 -422683
rect 34 -422717 46 -422683
rect -46 -422723 46 -422717
rect -102 -422767 -56 -422755
rect -102 -423743 -96 -422767
rect -62 -423743 -56 -422767
rect -102 -423755 -56 -423743
rect 56 -422767 102 -422755
rect 56 -423743 62 -422767
rect 96 -423743 102 -422767
rect 56 -423755 102 -423743
rect -46 -423793 46 -423787
rect -46 -423827 -34 -423793
rect 34 -423827 46 -423793
rect -46 -423833 46 -423827
rect -46 -423901 46 -423895
rect -46 -423935 -34 -423901
rect 34 -423935 46 -423901
rect -46 -423941 46 -423935
rect -102 -423985 -56 -423973
rect -102 -424961 -96 -423985
rect -62 -424961 -56 -423985
rect -102 -424973 -56 -424961
rect 56 -423985 102 -423973
rect 56 -424961 62 -423985
rect 96 -424961 102 -423985
rect 56 -424973 102 -424961
rect -46 -425011 46 -425005
rect -46 -425045 -34 -425011
rect 34 -425045 46 -425011
rect -46 -425051 46 -425045
rect -46 -425119 46 -425113
rect -46 -425153 -34 -425119
rect 34 -425153 46 -425119
rect -46 -425159 46 -425153
rect -102 -425203 -56 -425191
rect -102 -426179 -96 -425203
rect -62 -426179 -56 -425203
rect -102 -426191 -56 -426179
rect 56 -425203 102 -425191
rect 56 -426179 62 -425203
rect 96 -426179 102 -425203
rect 56 -426191 102 -426179
rect -46 -426229 46 -426223
rect -46 -426263 -34 -426229
rect 34 -426263 46 -426229
rect -46 -426269 46 -426263
rect -46 -426337 46 -426331
rect -46 -426371 -34 -426337
rect 34 -426371 46 -426337
rect -46 -426377 46 -426371
rect -102 -426421 -56 -426409
rect -102 -427397 -96 -426421
rect -62 -427397 -56 -426421
rect -102 -427409 -56 -427397
rect 56 -426421 102 -426409
rect 56 -427397 62 -426421
rect 96 -427397 102 -426421
rect 56 -427409 102 -427397
rect -46 -427447 46 -427441
rect -46 -427481 -34 -427447
rect 34 -427481 46 -427447
rect -46 -427487 46 -427481
rect -46 -427555 46 -427549
rect -46 -427589 -34 -427555
rect 34 -427589 46 -427555
rect -46 -427595 46 -427589
rect -102 -427639 -56 -427627
rect -102 -428615 -96 -427639
rect -62 -428615 -56 -427639
rect -102 -428627 -56 -428615
rect 56 -427639 102 -427627
rect 56 -428615 62 -427639
rect 96 -428615 102 -427639
rect 56 -428627 102 -428615
rect -46 -428665 46 -428659
rect -46 -428699 -34 -428665
rect 34 -428699 46 -428665
rect -46 -428705 46 -428699
rect -46 -428773 46 -428767
rect -46 -428807 -34 -428773
rect 34 -428807 46 -428773
rect -46 -428813 46 -428807
rect -102 -428857 -56 -428845
rect -102 -429833 -96 -428857
rect -62 -429833 -56 -428857
rect -102 -429845 -56 -429833
rect 56 -428857 102 -428845
rect 56 -429833 62 -428857
rect 96 -429833 102 -428857
rect 56 -429845 102 -429833
rect -46 -429883 46 -429877
rect -46 -429917 -34 -429883
rect 34 -429917 46 -429883
rect -46 -429923 46 -429917
rect -46 -429991 46 -429985
rect -46 -430025 -34 -429991
rect 34 -430025 46 -429991
rect -46 -430031 46 -430025
rect -102 -430075 -56 -430063
rect -102 -431051 -96 -430075
rect -62 -431051 -56 -430075
rect -102 -431063 -56 -431051
rect 56 -430075 102 -430063
rect 56 -431051 62 -430075
rect 96 -431051 102 -430075
rect 56 -431063 102 -431051
rect -46 -431101 46 -431095
rect -46 -431135 -34 -431101
rect 34 -431135 46 -431101
rect -46 -431141 46 -431135
rect -46 -431209 46 -431203
rect -46 -431243 -34 -431209
rect 34 -431243 46 -431209
rect -46 -431249 46 -431243
rect -102 -431293 -56 -431281
rect -102 -432269 -96 -431293
rect -62 -432269 -56 -431293
rect -102 -432281 -56 -432269
rect 56 -431293 102 -431281
rect 56 -432269 62 -431293
rect 96 -432269 102 -431293
rect 56 -432281 102 -432269
rect -46 -432319 46 -432313
rect -46 -432353 -34 -432319
rect 34 -432353 46 -432319
rect -46 -432359 46 -432353
rect -46 -432427 46 -432421
rect -46 -432461 -34 -432427
rect 34 -432461 46 -432427
rect -46 -432467 46 -432461
rect -102 -432511 -56 -432499
rect -102 -433487 -96 -432511
rect -62 -433487 -56 -432511
rect -102 -433499 -56 -433487
rect 56 -432511 102 -432499
rect 56 -433487 62 -432511
rect 96 -433487 102 -432511
rect 56 -433499 102 -433487
rect -46 -433537 46 -433531
rect -46 -433571 -34 -433537
rect 34 -433571 46 -433537
rect -46 -433577 46 -433571
rect -46 -433645 46 -433639
rect -46 -433679 -34 -433645
rect 34 -433679 46 -433645
rect -46 -433685 46 -433679
rect -102 -433729 -56 -433717
rect -102 -434705 -96 -433729
rect -62 -434705 -56 -433729
rect -102 -434717 -56 -434705
rect 56 -433729 102 -433717
rect 56 -434705 62 -433729
rect 96 -434705 102 -433729
rect 56 -434717 102 -434705
rect -46 -434755 46 -434749
rect -46 -434789 -34 -434755
rect 34 -434789 46 -434755
rect -46 -434795 46 -434789
rect -46 -434863 46 -434857
rect -46 -434897 -34 -434863
rect 34 -434897 46 -434863
rect -46 -434903 46 -434897
rect -102 -434947 -56 -434935
rect -102 -435923 -96 -434947
rect -62 -435923 -56 -434947
rect -102 -435935 -56 -435923
rect 56 -434947 102 -434935
rect 56 -435923 62 -434947
rect 96 -435923 102 -434947
rect 56 -435935 102 -435923
rect -46 -435973 46 -435967
rect -46 -436007 -34 -435973
rect 34 -436007 46 -435973
rect -46 -436013 46 -436007
rect -46 -436081 46 -436075
rect -46 -436115 -34 -436081
rect 34 -436115 46 -436081
rect -46 -436121 46 -436115
rect -102 -436165 -56 -436153
rect -102 -437141 -96 -436165
rect -62 -437141 -56 -436165
rect -102 -437153 -56 -437141
rect 56 -436165 102 -436153
rect 56 -437141 62 -436165
rect 96 -437141 102 -436165
rect 56 -437153 102 -437141
rect -46 -437191 46 -437185
rect -46 -437225 -34 -437191
rect 34 -437225 46 -437191
rect -46 -437231 46 -437225
rect -46 -437299 46 -437293
rect -46 -437333 -34 -437299
rect 34 -437333 46 -437299
rect -46 -437339 46 -437333
rect -102 -437383 -56 -437371
rect -102 -438359 -96 -437383
rect -62 -438359 -56 -437383
rect -102 -438371 -56 -438359
rect 56 -437383 102 -437371
rect 56 -438359 62 -437383
rect 96 -438359 102 -437383
rect 56 -438371 102 -438359
rect -46 -438409 46 -438403
rect -46 -438443 -34 -438409
rect 34 -438443 46 -438409
rect -46 -438449 46 -438443
rect -46 -438517 46 -438511
rect -46 -438551 -34 -438517
rect 34 -438551 46 -438517
rect -46 -438557 46 -438551
rect -102 -438601 -56 -438589
rect -102 -439577 -96 -438601
rect -62 -439577 -56 -438601
rect -102 -439589 -56 -439577
rect 56 -438601 102 -438589
rect 56 -439577 62 -438601
rect 96 -439577 102 -438601
rect 56 -439589 102 -439577
rect -46 -439627 46 -439621
rect -46 -439661 -34 -439627
rect 34 -439661 46 -439627
rect -46 -439667 46 -439661
rect -46 -439735 46 -439729
rect -46 -439769 -34 -439735
rect 34 -439769 46 -439735
rect -46 -439775 46 -439769
rect -102 -439819 -56 -439807
rect -102 -440795 -96 -439819
rect -62 -440795 -56 -439819
rect -102 -440807 -56 -440795
rect 56 -439819 102 -439807
rect 56 -440795 62 -439819
rect 96 -440795 102 -439819
rect 56 -440807 102 -440795
rect -46 -440845 46 -440839
rect -46 -440879 -34 -440845
rect 34 -440879 46 -440845
rect -46 -440885 46 -440879
rect -46 -440953 46 -440947
rect -46 -440987 -34 -440953
rect 34 -440987 46 -440953
rect -46 -440993 46 -440987
rect -102 -441037 -56 -441025
rect -102 -442013 -96 -441037
rect -62 -442013 -56 -441037
rect -102 -442025 -56 -442013
rect 56 -441037 102 -441025
rect 56 -442013 62 -441037
rect 96 -442013 102 -441037
rect 56 -442025 102 -442013
rect -46 -442063 46 -442057
rect -46 -442097 -34 -442063
rect 34 -442097 46 -442063
rect -46 -442103 46 -442097
rect -46 -442171 46 -442165
rect -46 -442205 -34 -442171
rect 34 -442205 46 -442171
rect -46 -442211 46 -442205
rect -102 -442255 -56 -442243
rect -102 -443231 -96 -442255
rect -62 -443231 -56 -442255
rect -102 -443243 -56 -443231
rect 56 -442255 102 -442243
rect 56 -443231 62 -442255
rect 96 -443231 102 -442255
rect 56 -443243 102 -443231
rect -46 -443281 46 -443275
rect -46 -443315 -34 -443281
rect 34 -443315 46 -443281
rect -46 -443321 46 -443315
rect -46 -443389 46 -443383
rect -46 -443423 -34 -443389
rect 34 -443423 46 -443389
rect -46 -443429 46 -443423
rect -102 -443473 -56 -443461
rect -102 -444449 -96 -443473
rect -62 -444449 -56 -443473
rect -102 -444461 -56 -444449
rect 56 -443473 102 -443461
rect 56 -444449 62 -443473
rect 96 -444449 102 -443473
rect 56 -444461 102 -444449
rect -46 -444499 46 -444493
rect -46 -444533 -34 -444499
rect 34 -444533 46 -444499
rect -46 -444539 46 -444533
rect -46 -444607 46 -444601
rect -46 -444641 -34 -444607
rect 34 -444641 46 -444607
rect -46 -444647 46 -444641
rect -102 -444691 -56 -444679
rect -102 -445667 -96 -444691
rect -62 -445667 -56 -444691
rect -102 -445679 -56 -445667
rect 56 -444691 102 -444679
rect 56 -445667 62 -444691
rect 96 -445667 102 -444691
rect 56 -445679 102 -445667
rect -46 -445717 46 -445711
rect -46 -445751 -34 -445717
rect 34 -445751 46 -445717
rect -46 -445757 46 -445751
rect -46 -445825 46 -445819
rect -46 -445859 -34 -445825
rect 34 -445859 46 -445825
rect -46 -445865 46 -445859
rect -102 -445909 -56 -445897
rect -102 -446885 -96 -445909
rect -62 -446885 -56 -445909
rect -102 -446897 -56 -446885
rect 56 -445909 102 -445897
rect 56 -446885 62 -445909
rect 96 -446885 102 -445909
rect 56 -446897 102 -446885
rect -46 -446935 46 -446929
rect -46 -446969 -34 -446935
rect 34 -446969 46 -446935
rect -46 -446975 46 -446969
rect -46 -447043 46 -447037
rect -46 -447077 -34 -447043
rect 34 -447077 46 -447043
rect -46 -447083 46 -447077
rect -102 -447127 -56 -447115
rect -102 -448103 -96 -447127
rect -62 -448103 -56 -447127
rect -102 -448115 -56 -448103
rect 56 -447127 102 -447115
rect 56 -448103 62 -447127
rect 96 -448103 102 -447127
rect 56 -448115 102 -448103
rect -46 -448153 46 -448147
rect -46 -448187 -34 -448153
rect 34 -448187 46 -448153
rect -46 -448193 46 -448187
rect -46 -448261 46 -448255
rect -46 -448295 -34 -448261
rect 34 -448295 46 -448261
rect -46 -448301 46 -448295
rect -102 -448345 -56 -448333
rect -102 -449321 -96 -448345
rect -62 -449321 -56 -448345
rect -102 -449333 -56 -449321
rect 56 -448345 102 -448333
rect 56 -449321 62 -448345
rect 96 -449321 102 -448345
rect 56 -449333 102 -449321
rect -46 -449371 46 -449365
rect -46 -449405 -34 -449371
rect 34 -449405 46 -449371
rect -46 -449411 46 -449405
rect -46 -449479 46 -449473
rect -46 -449513 -34 -449479
rect 34 -449513 46 -449479
rect -46 -449519 46 -449513
rect -102 -449563 -56 -449551
rect -102 -450539 -96 -449563
rect -62 -450539 -56 -449563
rect -102 -450551 -56 -450539
rect 56 -449563 102 -449551
rect 56 -450539 62 -449563
rect 96 -450539 102 -449563
rect 56 -450551 102 -450539
rect -46 -450589 46 -450583
rect -46 -450623 -34 -450589
rect 34 -450623 46 -450589
rect -46 -450629 46 -450623
rect -46 -450697 46 -450691
rect -46 -450731 -34 -450697
rect 34 -450731 46 -450697
rect -46 -450737 46 -450731
rect -102 -450781 -56 -450769
rect -102 -451757 -96 -450781
rect -62 -451757 -56 -450781
rect -102 -451769 -56 -451757
rect 56 -450781 102 -450769
rect 56 -451757 62 -450781
rect 96 -451757 102 -450781
rect 56 -451769 102 -451757
rect -46 -451807 46 -451801
rect -46 -451841 -34 -451807
rect 34 -451841 46 -451807
rect -46 -451847 46 -451841
rect -46 -451915 46 -451909
rect -46 -451949 -34 -451915
rect 34 -451949 46 -451915
rect -46 -451955 46 -451949
rect -102 -451999 -56 -451987
rect -102 -452975 -96 -451999
rect -62 -452975 -56 -451999
rect -102 -452987 -56 -452975
rect 56 -451999 102 -451987
rect 56 -452975 62 -451999
rect 96 -452975 102 -451999
rect 56 -452987 102 -452975
rect -46 -453025 46 -453019
rect -46 -453059 -34 -453025
rect 34 -453059 46 -453025
rect -46 -453065 46 -453059
rect -46 -453133 46 -453127
rect -46 -453167 -34 -453133
rect 34 -453167 46 -453133
rect -46 -453173 46 -453167
rect -102 -453217 -56 -453205
rect -102 -454193 -96 -453217
rect -62 -454193 -56 -453217
rect -102 -454205 -56 -454193
rect 56 -453217 102 -453205
rect 56 -454193 62 -453217
rect 96 -454193 102 -453217
rect 56 -454205 102 -454193
rect -46 -454243 46 -454237
rect -46 -454277 -34 -454243
rect 34 -454277 46 -454243
rect -46 -454283 46 -454277
rect -46 -454351 46 -454345
rect -46 -454385 -34 -454351
rect 34 -454385 46 -454351
rect -46 -454391 46 -454385
rect -102 -454435 -56 -454423
rect -102 -455411 -96 -454435
rect -62 -455411 -56 -454435
rect -102 -455423 -56 -455411
rect 56 -454435 102 -454423
rect 56 -455411 62 -454435
rect 96 -455411 102 -454435
rect 56 -455423 102 -455411
rect -46 -455461 46 -455455
rect -46 -455495 -34 -455461
rect 34 -455495 46 -455461
rect -46 -455501 46 -455495
rect -46 -455569 46 -455563
rect -46 -455603 -34 -455569
rect 34 -455603 46 -455569
rect -46 -455609 46 -455603
rect -102 -455653 -56 -455641
rect -102 -456629 -96 -455653
rect -62 -456629 -56 -455653
rect -102 -456641 -56 -456629
rect 56 -455653 102 -455641
rect 56 -456629 62 -455653
rect 96 -456629 102 -455653
rect 56 -456641 102 -456629
rect -46 -456679 46 -456673
rect -46 -456713 -34 -456679
rect 34 -456713 46 -456679
rect -46 -456719 46 -456713
rect -46 -456787 46 -456781
rect -46 -456821 -34 -456787
rect 34 -456821 46 -456787
rect -46 -456827 46 -456821
rect -102 -456871 -56 -456859
rect -102 -457847 -96 -456871
rect -62 -457847 -56 -456871
rect -102 -457859 -56 -457847
rect 56 -456871 102 -456859
rect 56 -457847 62 -456871
rect 96 -457847 102 -456871
rect 56 -457859 102 -457847
rect -46 -457897 46 -457891
rect -46 -457931 -34 -457897
rect 34 -457931 46 -457897
rect -46 -457937 46 -457931
rect -46 -458005 46 -457999
rect -46 -458039 -34 -458005
rect 34 -458039 46 -458005
rect -46 -458045 46 -458039
rect -102 -458089 -56 -458077
rect -102 -459065 -96 -458089
rect -62 -459065 -56 -458089
rect -102 -459077 -56 -459065
rect 56 -458089 102 -458077
rect 56 -459065 62 -458089
rect 96 -459065 102 -458089
rect 56 -459077 102 -459065
rect -46 -459115 46 -459109
rect -46 -459149 -34 -459115
rect 34 -459149 46 -459115
rect -46 -459155 46 -459149
rect -46 -459223 46 -459217
rect -46 -459257 -34 -459223
rect 34 -459257 46 -459223
rect -46 -459263 46 -459257
rect -102 -459307 -56 -459295
rect -102 -460283 -96 -459307
rect -62 -460283 -56 -459307
rect -102 -460295 -56 -460283
rect 56 -459307 102 -459295
rect 56 -460283 62 -459307
rect 96 -460283 102 -459307
rect 56 -460295 102 -460283
rect -46 -460333 46 -460327
rect -46 -460367 -34 -460333
rect 34 -460367 46 -460333
rect -46 -460373 46 -460367
rect -46 -460441 46 -460435
rect -46 -460475 -34 -460441
rect 34 -460475 46 -460441
rect -46 -460481 46 -460475
rect -102 -460525 -56 -460513
rect -102 -461501 -96 -460525
rect -62 -461501 -56 -460525
rect -102 -461513 -56 -461501
rect 56 -460525 102 -460513
rect 56 -461501 62 -460525
rect 96 -461501 102 -460525
rect 56 -461513 102 -461501
rect -46 -461551 46 -461545
rect -46 -461585 -34 -461551
rect 34 -461585 46 -461551
rect -46 -461591 46 -461585
rect -46 -461659 46 -461653
rect -46 -461693 -34 -461659
rect 34 -461693 46 -461659
rect -46 -461699 46 -461693
rect -102 -461743 -56 -461731
rect -102 -462719 -96 -461743
rect -62 -462719 -56 -461743
rect -102 -462731 -56 -462719
rect 56 -461743 102 -461731
rect 56 -462719 62 -461743
rect 96 -462719 102 -461743
rect 56 -462731 102 -462719
rect -46 -462769 46 -462763
rect -46 -462803 -34 -462769
rect 34 -462803 46 -462769
rect -46 -462809 46 -462803
rect -46 -462877 46 -462871
rect -46 -462911 -34 -462877
rect 34 -462911 46 -462877
rect -46 -462917 46 -462911
rect -102 -462961 -56 -462949
rect -102 -463937 -96 -462961
rect -62 -463937 -56 -462961
rect -102 -463949 -56 -463937
rect 56 -462961 102 -462949
rect 56 -463937 62 -462961
rect 96 -463937 102 -462961
rect 56 -463949 102 -463937
rect -46 -463987 46 -463981
rect -46 -464021 -34 -463987
rect 34 -464021 46 -463987
rect -46 -464027 46 -464021
rect -46 -464095 46 -464089
rect -46 -464129 -34 -464095
rect 34 -464129 46 -464095
rect -46 -464135 46 -464129
rect -102 -464179 -56 -464167
rect -102 -465155 -96 -464179
rect -62 -465155 -56 -464179
rect -102 -465167 -56 -465155
rect 56 -464179 102 -464167
rect 56 -465155 62 -464179
rect 96 -465155 102 -464179
rect 56 -465167 102 -465155
rect -46 -465205 46 -465199
rect -46 -465239 -34 -465205
rect 34 -465239 46 -465205
rect -46 -465245 46 -465239
rect -46 -465313 46 -465307
rect -46 -465347 -34 -465313
rect 34 -465347 46 -465313
rect -46 -465353 46 -465347
rect -102 -465397 -56 -465385
rect -102 -466373 -96 -465397
rect -62 -466373 -56 -465397
rect -102 -466385 -56 -466373
rect 56 -465397 102 -465385
rect 56 -466373 62 -465397
rect 96 -466373 102 -465397
rect 56 -466385 102 -466373
rect -46 -466423 46 -466417
rect -46 -466457 -34 -466423
rect 34 -466457 46 -466423
rect -46 -466463 46 -466457
rect -46 -466531 46 -466525
rect -46 -466565 -34 -466531
rect 34 -466565 46 -466531
rect -46 -466571 46 -466565
rect -102 -466615 -56 -466603
rect -102 -467591 -96 -466615
rect -62 -467591 -56 -466615
rect -102 -467603 -56 -467591
rect 56 -466615 102 -466603
rect 56 -467591 62 -466615
rect 96 -467591 102 -466615
rect 56 -467603 102 -467591
rect -46 -467641 46 -467635
rect -46 -467675 -34 -467641
rect 34 -467675 46 -467641
rect -46 -467681 46 -467675
rect -46 -467749 46 -467743
rect -46 -467783 -34 -467749
rect 34 -467783 46 -467749
rect -46 -467789 46 -467783
rect -102 -467833 -56 -467821
rect -102 -468809 -96 -467833
rect -62 -468809 -56 -467833
rect -102 -468821 -56 -468809
rect 56 -467833 102 -467821
rect 56 -468809 62 -467833
rect 96 -468809 102 -467833
rect 56 -468821 102 -468809
rect -46 -468859 46 -468853
rect -46 -468893 -34 -468859
rect 34 -468893 46 -468859
rect -46 -468899 46 -468893
rect -46 -468967 46 -468961
rect -46 -469001 -34 -468967
rect 34 -469001 46 -468967
rect -46 -469007 46 -469001
rect -102 -469051 -56 -469039
rect -102 -470027 -96 -469051
rect -62 -470027 -56 -469051
rect -102 -470039 -56 -470027
rect 56 -469051 102 -469039
rect 56 -470027 62 -469051
rect 96 -470027 102 -469051
rect 56 -470039 102 -470027
rect -46 -470077 46 -470071
rect -46 -470111 -34 -470077
rect 34 -470111 46 -470077
rect -46 -470117 46 -470111
rect -46 -470185 46 -470179
rect -46 -470219 -34 -470185
rect 34 -470219 46 -470185
rect -46 -470225 46 -470219
rect -102 -470269 -56 -470257
rect -102 -471245 -96 -470269
rect -62 -471245 -56 -470269
rect -102 -471257 -56 -471245
rect 56 -470269 102 -470257
rect 56 -471245 62 -470269
rect 96 -471245 102 -470269
rect 56 -471257 102 -471245
rect -46 -471295 46 -471289
rect -46 -471329 -34 -471295
rect 34 -471329 46 -471295
rect -46 -471335 46 -471329
rect -46 -471403 46 -471397
rect -46 -471437 -34 -471403
rect 34 -471437 46 -471403
rect -46 -471443 46 -471437
rect -102 -471487 -56 -471475
rect -102 -472463 -96 -471487
rect -62 -472463 -56 -471487
rect -102 -472475 -56 -472463
rect 56 -471487 102 -471475
rect 56 -472463 62 -471487
rect 96 -472463 102 -471487
rect 56 -472475 102 -472463
rect -46 -472513 46 -472507
rect -46 -472547 -34 -472513
rect 34 -472547 46 -472513
rect -46 -472553 46 -472547
rect -46 -472621 46 -472615
rect -46 -472655 -34 -472621
rect 34 -472655 46 -472621
rect -46 -472661 46 -472655
rect -102 -472705 -56 -472693
rect -102 -473681 -96 -472705
rect -62 -473681 -56 -472705
rect -102 -473693 -56 -473681
rect 56 -472705 102 -472693
rect 56 -473681 62 -472705
rect 96 -473681 102 -472705
rect 56 -473693 102 -473681
rect -46 -473731 46 -473725
rect -46 -473765 -34 -473731
rect 34 -473765 46 -473731
rect -46 -473771 46 -473765
rect -46 -473839 46 -473833
rect -46 -473873 -34 -473839
rect 34 -473873 46 -473839
rect -46 -473879 46 -473873
rect -102 -473923 -56 -473911
rect -102 -474899 -96 -473923
rect -62 -474899 -56 -473923
rect -102 -474911 -56 -474899
rect 56 -473923 102 -473911
rect 56 -474899 62 -473923
rect 96 -474899 102 -473923
rect 56 -474911 102 -474899
rect -46 -474949 46 -474943
rect -46 -474983 -34 -474949
rect 34 -474983 46 -474949
rect -46 -474989 46 -474983
rect -46 -475057 46 -475051
rect -46 -475091 -34 -475057
rect 34 -475091 46 -475057
rect -46 -475097 46 -475091
rect -102 -475141 -56 -475129
rect -102 -476117 -96 -475141
rect -62 -476117 -56 -475141
rect -102 -476129 -56 -476117
rect 56 -475141 102 -475129
rect 56 -476117 62 -475141
rect 96 -476117 102 -475141
rect 56 -476129 102 -476117
rect -46 -476167 46 -476161
rect -46 -476201 -34 -476167
rect 34 -476201 46 -476167
rect -46 -476207 46 -476201
rect -46 -476275 46 -476269
rect -46 -476309 -34 -476275
rect 34 -476309 46 -476275
rect -46 -476315 46 -476309
rect -102 -476359 -56 -476347
rect -102 -477335 -96 -476359
rect -62 -477335 -56 -476359
rect -102 -477347 -56 -477335
rect 56 -476359 102 -476347
rect 56 -477335 62 -476359
rect 96 -477335 102 -476359
rect 56 -477347 102 -477335
rect -46 -477385 46 -477379
rect -46 -477419 -34 -477385
rect 34 -477419 46 -477385
rect -46 -477425 46 -477419
rect -46 -477493 46 -477487
rect -46 -477527 -34 -477493
rect 34 -477527 46 -477493
rect -46 -477533 46 -477527
rect -102 -477577 -56 -477565
rect -102 -478553 -96 -477577
rect -62 -478553 -56 -477577
rect -102 -478565 -56 -478553
rect 56 -477577 102 -477565
rect 56 -478553 62 -477577
rect 96 -478553 102 -477577
rect 56 -478565 102 -478553
rect -46 -478603 46 -478597
rect -46 -478637 -34 -478603
rect 34 -478637 46 -478603
rect -46 -478643 46 -478637
rect -46 -478711 46 -478705
rect -46 -478745 -34 -478711
rect 34 -478745 46 -478711
rect -46 -478751 46 -478745
rect -102 -478795 -56 -478783
rect -102 -479771 -96 -478795
rect -62 -479771 -56 -478795
rect -102 -479783 -56 -479771
rect 56 -478795 102 -478783
rect 56 -479771 62 -478795
rect 96 -479771 102 -478795
rect 56 -479783 102 -479771
rect -46 -479821 46 -479815
rect -46 -479855 -34 -479821
rect 34 -479855 46 -479821
rect -46 -479861 46 -479855
rect -46 -479929 46 -479923
rect -46 -479963 -34 -479929
rect 34 -479963 46 -479929
rect -46 -479969 46 -479963
rect -102 -480013 -56 -480001
rect -102 -480989 -96 -480013
rect -62 -480989 -56 -480013
rect -102 -481001 -56 -480989
rect 56 -480013 102 -480001
rect 56 -480989 62 -480013
rect 96 -480989 102 -480013
rect 56 -481001 102 -480989
rect -46 -481039 46 -481033
rect -46 -481073 -34 -481039
rect 34 -481073 46 -481039
rect -46 -481079 46 -481073
rect -46 -481147 46 -481141
rect -46 -481181 -34 -481147
rect 34 -481181 46 -481147
rect -46 -481187 46 -481181
rect -102 -481231 -56 -481219
rect -102 -482207 -96 -481231
rect -62 -482207 -56 -481231
rect -102 -482219 -56 -482207
rect 56 -481231 102 -481219
rect 56 -482207 62 -481231
rect 96 -482207 102 -481231
rect 56 -482219 102 -482207
rect -46 -482257 46 -482251
rect -46 -482291 -34 -482257
rect 34 -482291 46 -482257
rect -46 -482297 46 -482291
rect -46 -482365 46 -482359
rect -46 -482399 -34 -482365
rect 34 -482399 46 -482365
rect -46 -482405 46 -482399
rect -102 -482449 -56 -482437
rect -102 -483425 -96 -482449
rect -62 -483425 -56 -482449
rect -102 -483437 -56 -483425
rect 56 -482449 102 -482437
rect 56 -483425 62 -482449
rect 96 -483425 102 -482449
rect 56 -483437 102 -483425
rect -46 -483475 46 -483469
rect -46 -483509 -34 -483475
rect 34 -483509 46 -483475
rect -46 -483515 46 -483509
rect -46 -483583 46 -483577
rect -46 -483617 -34 -483583
rect 34 -483617 46 -483583
rect -46 -483623 46 -483617
rect -102 -483667 -56 -483655
rect -102 -484643 -96 -483667
rect -62 -484643 -56 -483667
rect -102 -484655 -56 -484643
rect 56 -483667 102 -483655
rect 56 -484643 62 -483667
rect 96 -484643 102 -483667
rect 56 -484655 102 -484643
rect -46 -484693 46 -484687
rect -46 -484727 -34 -484693
rect 34 -484727 46 -484693
rect -46 -484733 46 -484727
rect -46 -484801 46 -484795
rect -46 -484835 -34 -484801
rect 34 -484835 46 -484801
rect -46 -484841 46 -484835
rect -102 -484885 -56 -484873
rect -102 -485861 -96 -484885
rect -62 -485861 -56 -484885
rect -102 -485873 -56 -485861
rect 56 -484885 102 -484873
rect 56 -485861 62 -484885
rect 96 -485861 102 -484885
rect 56 -485873 102 -485861
rect -46 -485911 46 -485905
rect -46 -485945 -34 -485911
rect 34 -485945 46 -485911
rect -46 -485951 46 -485945
rect -46 -486019 46 -486013
rect -46 -486053 -34 -486019
rect 34 -486053 46 -486019
rect -46 -486059 46 -486053
rect -102 -486103 -56 -486091
rect -102 -487079 -96 -486103
rect -62 -487079 -56 -486103
rect -102 -487091 -56 -487079
rect 56 -486103 102 -486091
rect 56 -487079 62 -486103
rect 96 -487079 102 -486103
rect 56 -487091 102 -487079
rect -46 -487129 46 -487123
rect -46 -487163 -34 -487129
rect 34 -487163 46 -487129
rect -46 -487169 46 -487163
rect -46 -487237 46 -487231
rect -46 -487271 -34 -487237
rect 34 -487271 46 -487237
rect -46 -487277 46 -487271
rect -102 -487321 -56 -487309
rect -102 -488297 -96 -487321
rect -62 -488297 -56 -487321
rect -102 -488309 -56 -488297
rect 56 -487321 102 -487309
rect 56 -488297 62 -487321
rect 96 -488297 102 -487321
rect 56 -488309 102 -488297
rect -46 -488347 46 -488341
rect -46 -488381 -34 -488347
rect 34 -488381 46 -488347
rect -46 -488387 46 -488381
rect -46 -488455 46 -488449
rect -46 -488489 -34 -488455
rect 34 -488489 46 -488455
rect -46 -488495 46 -488489
rect -102 -488539 -56 -488527
rect -102 -489515 -96 -488539
rect -62 -489515 -56 -488539
rect -102 -489527 -56 -489515
rect 56 -488539 102 -488527
rect 56 -489515 62 -488539
rect 96 -489515 102 -488539
rect 56 -489527 102 -489515
rect -46 -489565 46 -489559
rect -46 -489599 -34 -489565
rect 34 -489599 46 -489565
rect -46 -489605 46 -489599
rect -46 -489673 46 -489667
rect -46 -489707 -34 -489673
rect 34 -489707 46 -489673
rect -46 -489713 46 -489707
rect -102 -489757 -56 -489745
rect -102 -490733 -96 -489757
rect -62 -490733 -56 -489757
rect -102 -490745 -56 -490733
rect 56 -489757 102 -489745
rect 56 -490733 62 -489757
rect 96 -490733 102 -489757
rect 56 -490745 102 -490733
rect -46 -490783 46 -490777
rect -46 -490817 -34 -490783
rect 34 -490817 46 -490783
rect -46 -490823 46 -490817
rect -46 -490891 46 -490885
rect -46 -490925 -34 -490891
rect 34 -490925 46 -490891
rect -46 -490931 46 -490925
rect -102 -490975 -56 -490963
rect -102 -491951 -96 -490975
rect -62 -491951 -56 -490975
rect -102 -491963 -56 -491951
rect 56 -490975 102 -490963
rect 56 -491951 62 -490975
rect 96 -491951 102 -490975
rect 56 -491963 102 -491951
rect -46 -492001 46 -491995
rect -46 -492035 -34 -492001
rect 34 -492035 46 -492001
rect -46 -492041 46 -492035
rect -46 -492109 46 -492103
rect -46 -492143 -34 -492109
rect 34 -492143 46 -492109
rect -46 -492149 46 -492143
rect -102 -492193 -56 -492181
rect -102 -493169 -96 -492193
rect -62 -493169 -56 -492193
rect -102 -493181 -56 -493169
rect 56 -492193 102 -492181
rect 56 -493169 62 -492193
rect 96 -493169 102 -492193
rect 56 -493181 102 -493169
rect -46 -493219 46 -493213
rect -46 -493253 -34 -493219
rect 34 -493253 46 -493219
rect -46 -493259 46 -493253
rect -46 -493327 46 -493321
rect -46 -493361 -34 -493327
rect 34 -493361 46 -493327
rect -46 -493367 46 -493361
rect -102 -493411 -56 -493399
rect -102 -494387 -96 -493411
rect -62 -494387 -56 -493411
rect -102 -494399 -56 -494387
rect 56 -493411 102 -493399
rect 56 -494387 62 -493411
rect 96 -494387 102 -493411
rect 56 -494399 102 -494387
rect -46 -494437 46 -494431
rect -46 -494471 -34 -494437
rect 34 -494471 46 -494437
rect -46 -494477 46 -494471
rect -46 -494545 46 -494539
rect -46 -494579 -34 -494545
rect 34 -494579 46 -494545
rect -46 -494585 46 -494579
rect -102 -494629 -56 -494617
rect -102 -495605 -96 -494629
rect -62 -495605 -56 -494629
rect -102 -495617 -56 -495605
rect 56 -494629 102 -494617
rect 56 -495605 62 -494629
rect 96 -495605 102 -494629
rect 56 -495617 102 -495605
rect -46 -495655 46 -495649
rect -46 -495689 -34 -495655
rect 34 -495689 46 -495655
rect -46 -495695 46 -495689
rect -46 -495763 46 -495757
rect -46 -495797 -34 -495763
rect 34 -495797 46 -495763
rect -46 -495803 46 -495797
rect -102 -495847 -56 -495835
rect -102 -496823 -96 -495847
rect -62 -496823 -56 -495847
rect -102 -496835 -56 -496823
rect 56 -495847 102 -495835
rect 56 -496823 62 -495847
rect 96 -496823 102 -495847
rect 56 -496835 102 -496823
rect -46 -496873 46 -496867
rect -46 -496907 -34 -496873
rect 34 -496907 46 -496873
rect -46 -496913 46 -496907
rect -46 -496981 46 -496975
rect -46 -497015 -34 -496981
rect 34 -497015 46 -496981
rect -46 -497021 46 -497015
rect -102 -497065 -56 -497053
rect -102 -498041 -96 -497065
rect -62 -498041 -56 -497065
rect -102 -498053 -56 -498041
rect 56 -497065 102 -497053
rect 56 -498041 62 -497065
rect 96 -498041 102 -497065
rect 56 -498053 102 -498041
rect -46 -498091 46 -498085
rect -46 -498125 -34 -498091
rect 34 -498125 46 -498091
rect -46 -498131 46 -498125
rect -46 -498199 46 -498193
rect -46 -498233 -34 -498199
rect 34 -498233 46 -498199
rect -46 -498239 46 -498233
rect -102 -498283 -56 -498271
rect -102 -499259 -96 -498283
rect -62 -499259 -56 -498283
rect -102 -499271 -56 -499259
rect 56 -498283 102 -498271
rect 56 -499259 62 -498283
rect 96 -499259 102 -498283
rect 56 -499271 102 -499259
rect -46 -499309 46 -499303
rect -46 -499343 -34 -499309
rect 34 -499343 46 -499309
rect -46 -499349 46 -499343
rect -46 -499417 46 -499411
rect -46 -499451 -34 -499417
rect 34 -499451 46 -499417
rect -46 -499457 46 -499451
rect -102 -499501 -56 -499489
rect -102 -500477 -96 -499501
rect -62 -500477 -56 -499501
rect -102 -500489 -56 -500477
rect 56 -499501 102 -499489
rect 56 -500477 62 -499501
rect 96 -500477 102 -499501
rect 56 -500489 102 -500477
rect -46 -500527 46 -500521
rect -46 -500561 -34 -500527
rect 34 -500561 46 -500527
rect -46 -500567 46 -500561
rect -46 -500635 46 -500629
rect -46 -500669 -34 -500635
rect 34 -500669 46 -500635
rect -46 -500675 46 -500669
rect -102 -500719 -56 -500707
rect -102 -501695 -96 -500719
rect -62 -501695 -56 -500719
rect -102 -501707 -56 -501695
rect 56 -500719 102 -500707
rect 56 -501695 62 -500719
rect 96 -501695 102 -500719
rect 56 -501707 102 -501695
rect -46 -501745 46 -501739
rect -46 -501779 -34 -501745
rect 34 -501779 46 -501745
rect -46 -501785 46 -501779
rect -46 -501853 46 -501847
rect -46 -501887 -34 -501853
rect 34 -501887 46 -501853
rect -46 -501893 46 -501887
rect -102 -501937 -56 -501925
rect -102 -502913 -96 -501937
rect -62 -502913 -56 -501937
rect -102 -502925 -56 -502913
rect 56 -501937 102 -501925
rect 56 -502913 62 -501937
rect 96 -502913 102 -501937
rect 56 -502925 102 -502913
rect -46 -502963 46 -502957
rect -46 -502997 -34 -502963
rect 34 -502997 46 -502963
rect -46 -503003 46 -502997
rect -46 -503071 46 -503065
rect -46 -503105 -34 -503071
rect 34 -503105 46 -503071
rect -46 -503111 46 -503105
rect -102 -503155 -56 -503143
rect -102 -504131 -96 -503155
rect -62 -504131 -56 -503155
rect -102 -504143 -56 -504131
rect 56 -503155 102 -503143
rect 56 -504131 62 -503155
rect 96 -504131 102 -503155
rect 56 -504143 102 -504131
rect -46 -504181 46 -504175
rect -46 -504215 -34 -504181
rect 34 -504215 46 -504181
rect -46 -504221 46 -504215
rect -46 -504289 46 -504283
rect -46 -504323 -34 -504289
rect 34 -504323 46 -504289
rect -46 -504329 46 -504323
rect -102 -504373 -56 -504361
rect -102 -505349 -96 -504373
rect -62 -505349 -56 -504373
rect -102 -505361 -56 -505349
rect 56 -504373 102 -504361
rect 56 -505349 62 -504373
rect 96 -505349 102 -504373
rect 56 -505361 102 -505349
rect -46 -505399 46 -505393
rect -46 -505433 -34 -505399
rect 34 -505433 46 -505399
rect -46 -505439 46 -505433
rect -46 -505507 46 -505501
rect -46 -505541 -34 -505507
rect 34 -505541 46 -505507
rect -46 -505547 46 -505541
rect -102 -505591 -56 -505579
rect -102 -506567 -96 -505591
rect -62 -506567 -56 -505591
rect -102 -506579 -56 -506567
rect 56 -505591 102 -505579
rect 56 -506567 62 -505591
rect 96 -506567 102 -505591
rect 56 -506579 102 -506567
rect -46 -506617 46 -506611
rect -46 -506651 -34 -506617
rect 34 -506651 46 -506617
rect -46 -506657 46 -506651
rect -46 -506725 46 -506719
rect -46 -506759 -34 -506725
rect 34 -506759 46 -506725
rect -46 -506765 46 -506759
rect -102 -506809 -56 -506797
rect -102 -507785 -96 -506809
rect -62 -507785 -56 -506809
rect -102 -507797 -56 -507785
rect 56 -506809 102 -506797
rect 56 -507785 62 -506809
rect 96 -507785 102 -506809
rect 56 -507797 102 -507785
rect -46 -507835 46 -507829
rect -46 -507869 -34 -507835
rect 34 -507869 46 -507835
rect -46 -507875 46 -507869
rect -46 -507943 46 -507937
rect -46 -507977 -34 -507943
rect 34 -507977 46 -507943
rect -46 -507983 46 -507977
rect -102 -508027 -56 -508015
rect -102 -509003 -96 -508027
rect -62 -509003 -56 -508027
rect -102 -509015 -56 -509003
rect 56 -508027 102 -508015
rect 56 -509003 62 -508027
rect 96 -509003 102 -508027
rect 56 -509015 102 -509003
rect -46 -509053 46 -509047
rect -46 -509087 -34 -509053
rect 34 -509087 46 -509053
rect -46 -509093 46 -509087
rect -46 -509161 46 -509155
rect -46 -509195 -34 -509161
rect 34 -509195 46 -509161
rect -46 -509201 46 -509195
rect -102 -509245 -56 -509233
rect -102 -510221 -96 -509245
rect -62 -510221 -56 -509245
rect -102 -510233 -56 -510221
rect 56 -509245 102 -509233
rect 56 -510221 62 -509245
rect 96 -510221 102 -509245
rect 56 -510233 102 -510221
rect -46 -510271 46 -510265
rect -46 -510305 -34 -510271
rect 34 -510305 46 -510271
rect -46 -510311 46 -510305
rect -46 -510379 46 -510373
rect -46 -510413 -34 -510379
rect 34 -510413 46 -510379
rect -46 -510419 46 -510413
rect -102 -510463 -56 -510451
rect -102 -511439 -96 -510463
rect -62 -511439 -56 -510463
rect -102 -511451 -56 -511439
rect 56 -510463 102 -510451
rect 56 -511439 62 -510463
rect 96 -511439 102 -510463
rect 56 -511451 102 -511439
rect -46 -511489 46 -511483
rect -46 -511523 -34 -511489
rect 34 -511523 46 -511489
rect -46 -511529 46 -511523
rect -46 -511597 46 -511591
rect -46 -511631 -34 -511597
rect 34 -511631 46 -511597
rect -46 -511637 46 -511631
rect -102 -511681 -56 -511669
rect -102 -512657 -96 -511681
rect -62 -512657 -56 -511681
rect -102 -512669 -56 -512657
rect 56 -511681 102 -511669
rect 56 -512657 62 -511681
rect 96 -512657 102 -511681
rect 56 -512669 102 -512657
rect -46 -512707 46 -512701
rect -46 -512741 -34 -512707
rect 34 -512741 46 -512707
rect -46 -512747 46 -512741
rect -46 -512815 46 -512809
rect -46 -512849 -34 -512815
rect 34 -512849 46 -512815
rect -46 -512855 46 -512849
rect -102 -512899 -56 -512887
rect -102 -513875 -96 -512899
rect -62 -513875 -56 -512899
rect -102 -513887 -56 -513875
rect 56 -512899 102 -512887
rect 56 -513875 62 -512899
rect 96 -513875 102 -512899
rect 56 -513887 102 -513875
rect -46 -513925 46 -513919
rect -46 -513959 -34 -513925
rect 34 -513959 46 -513925
rect -46 -513965 46 -513959
rect -46 -514033 46 -514027
rect -46 -514067 -34 -514033
rect 34 -514067 46 -514033
rect -46 -514073 46 -514067
rect -102 -514117 -56 -514105
rect -102 -515093 -96 -514117
rect -62 -515093 -56 -514117
rect -102 -515105 -56 -515093
rect 56 -514117 102 -514105
rect 56 -515093 62 -514117
rect 96 -515093 102 -514117
rect 56 -515105 102 -515093
rect -46 -515143 46 -515137
rect -46 -515177 -34 -515143
rect 34 -515177 46 -515143
rect -46 -515183 46 -515177
rect -46 -515251 46 -515245
rect -46 -515285 -34 -515251
rect 34 -515285 46 -515251
rect -46 -515291 46 -515285
rect -102 -515335 -56 -515323
rect -102 -516311 -96 -515335
rect -62 -516311 -56 -515335
rect -102 -516323 -56 -516311
rect 56 -515335 102 -515323
rect 56 -516311 62 -515335
rect 96 -516311 102 -515335
rect 56 -516323 102 -516311
rect -46 -516361 46 -516355
rect -46 -516395 -34 -516361
rect 34 -516395 46 -516361
rect -46 -516401 46 -516395
rect -46 -516469 46 -516463
rect -46 -516503 -34 -516469
rect 34 -516503 46 -516469
rect -46 -516509 46 -516503
rect -102 -516553 -56 -516541
rect -102 -517529 -96 -516553
rect -62 -517529 -56 -516553
rect -102 -517541 -56 -517529
rect 56 -516553 102 -516541
rect 56 -517529 62 -516553
rect 96 -517529 102 -516553
rect 56 -517541 102 -517529
rect -46 -517579 46 -517573
rect -46 -517613 -34 -517579
rect 34 -517613 46 -517579
rect -46 -517619 46 -517613
rect -46 -517687 46 -517681
rect -46 -517721 -34 -517687
rect 34 -517721 46 -517687
rect -46 -517727 46 -517721
rect -102 -517771 -56 -517759
rect -102 -518747 -96 -517771
rect -62 -518747 -56 -517771
rect -102 -518759 -56 -518747
rect 56 -517771 102 -517759
rect 56 -518747 62 -517771
rect 96 -518747 102 -517771
rect 56 -518759 102 -518747
rect -46 -518797 46 -518791
rect -46 -518831 -34 -518797
rect 34 -518831 46 -518797
rect -46 -518837 46 -518831
rect -46 -518905 46 -518899
rect -46 -518939 -34 -518905
rect 34 -518939 46 -518905
rect -46 -518945 46 -518939
rect -102 -518989 -56 -518977
rect -102 -519965 -96 -518989
rect -62 -519965 -56 -518989
rect -102 -519977 -56 -519965
rect 56 -518989 102 -518977
rect 56 -519965 62 -518989
rect 96 -519965 102 -518989
rect 56 -519977 102 -519965
rect -46 -520015 46 -520009
rect -46 -520049 -34 -520015
rect 34 -520049 46 -520015
rect -46 -520055 46 -520049
rect -46 -520123 46 -520117
rect -46 -520157 -34 -520123
rect 34 -520157 46 -520123
rect -46 -520163 46 -520157
rect -102 -520207 -56 -520195
rect -102 -521183 -96 -520207
rect -62 -521183 -56 -520207
rect -102 -521195 -56 -521183
rect 56 -520207 102 -520195
rect 56 -521183 62 -520207
rect 96 -521183 102 -520207
rect 56 -521195 102 -521183
rect -46 -521233 46 -521227
rect -46 -521267 -34 -521233
rect 34 -521267 46 -521233
rect -46 -521273 46 -521267
rect -46 -521341 46 -521335
rect -46 -521375 -34 -521341
rect 34 -521375 46 -521341
rect -46 -521381 46 -521375
rect -102 -521425 -56 -521413
rect -102 -522401 -96 -521425
rect -62 -522401 -56 -521425
rect -102 -522413 -56 -522401
rect 56 -521425 102 -521413
rect 56 -522401 62 -521425
rect 96 -522401 102 -521425
rect 56 -522413 102 -522401
rect -46 -522451 46 -522445
rect -46 -522485 -34 -522451
rect 34 -522485 46 -522451
rect -46 -522491 46 -522485
rect -46 -522559 46 -522553
rect -46 -522593 -34 -522559
rect 34 -522593 46 -522559
rect -46 -522599 46 -522593
rect -102 -522643 -56 -522631
rect -102 -523619 -96 -522643
rect -62 -523619 -56 -522643
rect -102 -523631 -56 -523619
rect 56 -522643 102 -522631
rect 56 -523619 62 -522643
rect 96 -523619 102 -522643
rect 56 -523631 102 -523619
rect -46 -523669 46 -523663
rect -46 -523703 -34 -523669
rect 34 -523703 46 -523669
rect -46 -523709 46 -523703
rect -46 -523777 46 -523771
rect -46 -523811 -34 -523777
rect 34 -523811 46 -523777
rect -46 -523817 46 -523811
rect -102 -523861 -56 -523849
rect -102 -524837 -96 -523861
rect -62 -524837 -56 -523861
rect -102 -524849 -56 -524837
rect 56 -523861 102 -523849
rect 56 -524837 62 -523861
rect 96 -524837 102 -523861
rect 56 -524849 102 -524837
rect -46 -524887 46 -524881
rect -46 -524921 -34 -524887
rect 34 -524921 46 -524887
rect -46 -524927 46 -524921
rect -46 -524995 46 -524989
rect -46 -525029 -34 -524995
rect 34 -525029 46 -524995
rect -46 -525035 46 -525029
rect -102 -525079 -56 -525067
rect -102 -526055 -96 -525079
rect -62 -526055 -56 -525079
rect -102 -526067 -56 -526055
rect 56 -525079 102 -525067
rect 56 -526055 62 -525079
rect 96 -526055 102 -525079
rect 56 -526067 102 -526055
rect -46 -526105 46 -526099
rect -46 -526139 -34 -526105
rect 34 -526139 46 -526105
rect -46 -526145 46 -526139
rect -46 -526213 46 -526207
rect -46 -526247 -34 -526213
rect 34 -526247 46 -526213
rect -46 -526253 46 -526247
rect -102 -526297 -56 -526285
rect -102 -527273 -96 -526297
rect -62 -527273 -56 -526297
rect -102 -527285 -56 -527273
rect 56 -526297 102 -526285
rect 56 -527273 62 -526297
rect 96 -527273 102 -526297
rect 56 -527285 102 -527273
rect -46 -527323 46 -527317
rect -46 -527357 -34 -527323
rect 34 -527357 46 -527323
rect -46 -527363 46 -527357
rect -46 -527431 46 -527425
rect -46 -527465 -34 -527431
rect 34 -527465 46 -527431
rect -46 -527471 46 -527465
rect -102 -527515 -56 -527503
rect -102 -528491 -96 -527515
rect -62 -528491 -56 -527515
rect -102 -528503 -56 -528491
rect 56 -527515 102 -527503
rect 56 -528491 62 -527515
rect 96 -528491 102 -527515
rect 56 -528503 102 -528491
rect -46 -528541 46 -528535
rect -46 -528575 -34 -528541
rect 34 -528575 46 -528541
rect -46 -528581 46 -528575
rect -46 -528649 46 -528643
rect -46 -528683 -34 -528649
rect 34 -528683 46 -528649
rect -46 -528689 46 -528683
rect -102 -528733 -56 -528721
rect -102 -529709 -96 -528733
rect -62 -529709 -56 -528733
rect -102 -529721 -56 -529709
rect 56 -528733 102 -528721
rect 56 -529709 62 -528733
rect 96 -529709 102 -528733
rect 56 -529721 102 -529709
rect -46 -529759 46 -529753
rect -46 -529793 -34 -529759
rect 34 -529793 46 -529759
rect -46 -529799 46 -529793
rect -46 -529867 46 -529861
rect -46 -529901 -34 -529867
rect 34 -529901 46 -529867
rect -46 -529907 46 -529901
rect -102 -529951 -56 -529939
rect -102 -530927 -96 -529951
rect -62 -530927 -56 -529951
rect -102 -530939 -56 -530927
rect 56 -529951 102 -529939
rect 56 -530927 62 -529951
rect 96 -530927 102 -529951
rect 56 -530939 102 -530927
rect -46 -530977 46 -530971
rect -46 -531011 -34 -530977
rect 34 -531011 46 -530977
rect -46 -531017 46 -531011
rect -46 -531085 46 -531079
rect -46 -531119 -34 -531085
rect 34 -531119 46 -531085
rect -46 -531125 46 -531119
rect -102 -531169 -56 -531157
rect -102 -532145 -96 -531169
rect -62 -532145 -56 -531169
rect -102 -532157 -56 -532145
rect 56 -531169 102 -531157
rect 56 -532145 62 -531169
rect 96 -532145 102 -531169
rect 56 -532157 102 -532145
rect -46 -532195 46 -532189
rect -46 -532229 -34 -532195
rect 34 -532229 46 -532195
rect -46 -532235 46 -532229
rect -46 -532303 46 -532297
rect -46 -532337 -34 -532303
rect 34 -532337 46 -532303
rect -46 -532343 46 -532337
rect -102 -532387 -56 -532375
rect -102 -533363 -96 -532387
rect -62 -533363 -56 -532387
rect -102 -533375 -56 -533363
rect 56 -532387 102 -532375
rect 56 -533363 62 -532387
rect 96 -533363 102 -532387
rect 56 -533375 102 -533363
rect -46 -533413 46 -533407
rect -46 -533447 -34 -533413
rect 34 -533447 46 -533413
rect -46 -533453 46 -533447
rect -46 -533521 46 -533515
rect -46 -533555 -34 -533521
rect 34 -533555 46 -533521
rect -46 -533561 46 -533555
rect -102 -533605 -56 -533593
rect -102 -534581 -96 -533605
rect -62 -534581 -56 -533605
rect -102 -534593 -56 -534581
rect 56 -533605 102 -533593
rect 56 -534581 62 -533605
rect 96 -534581 102 -533605
rect 56 -534593 102 -534581
rect -46 -534631 46 -534625
rect -46 -534665 -34 -534631
rect 34 -534665 46 -534631
rect -46 -534671 46 -534665
rect -46 -534739 46 -534733
rect -46 -534773 -34 -534739
rect 34 -534773 46 -534739
rect -46 -534779 46 -534773
rect -102 -534823 -56 -534811
rect -102 -535799 -96 -534823
rect -62 -535799 -56 -534823
rect -102 -535811 -56 -535799
rect 56 -534823 102 -534811
rect 56 -535799 62 -534823
rect 96 -535799 102 -534823
rect 56 -535811 102 -535799
rect -46 -535849 46 -535843
rect -46 -535883 -34 -535849
rect 34 -535883 46 -535849
rect -46 -535889 46 -535883
rect -46 -535957 46 -535951
rect -46 -535991 -34 -535957
rect 34 -535991 46 -535957
rect -46 -535997 46 -535991
rect -102 -536041 -56 -536029
rect -102 -537017 -96 -536041
rect -62 -537017 -56 -536041
rect -102 -537029 -56 -537017
rect 56 -536041 102 -536029
rect 56 -537017 62 -536041
rect 96 -537017 102 -536041
rect 56 -537029 102 -537017
rect -46 -537067 46 -537061
rect -46 -537101 -34 -537067
rect 34 -537101 46 -537067
rect -46 -537107 46 -537101
rect -46 -537175 46 -537169
rect -46 -537209 -34 -537175
rect 34 -537209 46 -537175
rect -46 -537215 46 -537209
rect -102 -537259 -56 -537247
rect -102 -538235 -96 -537259
rect -62 -538235 -56 -537259
rect -102 -538247 -56 -538235
rect 56 -537259 102 -537247
rect 56 -538235 62 -537259
rect 96 -538235 102 -537259
rect 56 -538247 102 -538235
rect -46 -538285 46 -538279
rect -46 -538319 -34 -538285
rect 34 -538319 46 -538285
rect -46 -538325 46 -538319
rect -46 -538393 46 -538387
rect -46 -538427 -34 -538393
rect 34 -538427 46 -538393
rect -46 -538433 46 -538427
rect -102 -538477 -56 -538465
rect -102 -539453 -96 -538477
rect -62 -539453 -56 -538477
rect -102 -539465 -56 -539453
rect 56 -538477 102 -538465
rect 56 -539453 62 -538477
rect 96 -539453 102 -538477
rect 56 -539465 102 -539453
rect -46 -539503 46 -539497
rect -46 -539537 -34 -539503
rect 34 -539537 46 -539503
rect -46 -539543 46 -539537
rect -46 -539611 46 -539605
rect -46 -539645 -34 -539611
rect 34 -539645 46 -539611
rect -46 -539651 46 -539645
rect -102 -539695 -56 -539683
rect -102 -540671 -96 -539695
rect -62 -540671 -56 -539695
rect -102 -540683 -56 -540671
rect 56 -539695 102 -539683
rect 56 -540671 62 -539695
rect 96 -540671 102 -539695
rect 56 -540683 102 -540671
rect -46 -540721 46 -540715
rect -46 -540755 -34 -540721
rect 34 -540755 46 -540721
rect -46 -540761 46 -540755
rect -46 -540829 46 -540823
rect -46 -540863 -34 -540829
rect 34 -540863 46 -540829
rect -46 -540869 46 -540863
rect -102 -540913 -56 -540901
rect -102 -541889 -96 -540913
rect -62 -541889 -56 -540913
rect -102 -541901 -56 -541889
rect 56 -540913 102 -540901
rect 56 -541889 62 -540913
rect 96 -541889 102 -540913
rect 56 -541901 102 -541889
rect -46 -541939 46 -541933
rect -46 -541973 -34 -541939
rect 34 -541973 46 -541939
rect -46 -541979 46 -541973
rect -46 -542047 46 -542041
rect -46 -542081 -34 -542047
rect 34 -542081 46 -542047
rect -46 -542087 46 -542081
rect -102 -542131 -56 -542119
rect -102 -543107 -96 -542131
rect -62 -543107 -56 -542131
rect -102 -543119 -56 -543107
rect 56 -542131 102 -542119
rect 56 -543107 62 -542131
rect 96 -543107 102 -542131
rect 56 -543119 102 -543107
rect -46 -543157 46 -543151
rect -46 -543191 -34 -543157
rect 34 -543191 46 -543157
rect -46 -543197 46 -543191
rect -46 -543265 46 -543259
rect -46 -543299 -34 -543265
rect 34 -543299 46 -543265
rect -46 -543305 46 -543299
rect -102 -543349 -56 -543337
rect -102 -544325 -96 -543349
rect -62 -544325 -56 -543349
rect -102 -544337 -56 -544325
rect 56 -543349 102 -543337
rect 56 -544325 62 -543349
rect 96 -544325 102 -543349
rect 56 -544337 102 -544325
rect -46 -544375 46 -544369
rect -46 -544409 -34 -544375
rect 34 -544409 46 -544375
rect -46 -544415 46 -544409
rect -46 -544483 46 -544477
rect -46 -544517 -34 -544483
rect 34 -544517 46 -544483
rect -46 -544523 46 -544517
rect -102 -544567 -56 -544555
rect -102 -545543 -96 -544567
rect -62 -545543 -56 -544567
rect -102 -545555 -56 -545543
rect 56 -544567 102 -544555
rect 56 -545543 62 -544567
rect 96 -545543 102 -544567
rect 56 -545555 102 -545543
rect -46 -545593 46 -545587
rect -46 -545627 -34 -545593
rect 34 -545627 46 -545593
rect -46 -545633 46 -545627
rect -46 -545701 46 -545695
rect -46 -545735 -34 -545701
rect 34 -545735 46 -545701
rect -46 -545741 46 -545735
rect -102 -545785 -56 -545773
rect -102 -546761 -96 -545785
rect -62 -546761 -56 -545785
rect -102 -546773 -56 -546761
rect 56 -545785 102 -545773
rect 56 -546761 62 -545785
rect 96 -546761 102 -545785
rect 56 -546773 102 -546761
rect -46 -546811 46 -546805
rect -46 -546845 -34 -546811
rect 34 -546845 46 -546811
rect -46 -546851 46 -546845
rect -46 -546919 46 -546913
rect -46 -546953 -34 -546919
rect 34 -546953 46 -546919
rect -46 -546959 46 -546953
rect -102 -547003 -56 -546991
rect -102 -547979 -96 -547003
rect -62 -547979 -56 -547003
rect -102 -547991 -56 -547979
rect 56 -547003 102 -546991
rect 56 -547979 62 -547003
rect 96 -547979 102 -547003
rect 56 -547991 102 -547979
rect -46 -548029 46 -548023
rect -46 -548063 -34 -548029
rect 34 -548063 46 -548029
rect -46 -548069 46 -548063
rect -46 -548137 46 -548131
rect -46 -548171 -34 -548137
rect 34 -548171 46 -548137
rect -46 -548177 46 -548171
rect -102 -548221 -56 -548209
rect -102 -549197 -96 -548221
rect -62 -549197 -56 -548221
rect -102 -549209 -56 -549197
rect 56 -548221 102 -548209
rect 56 -549197 62 -548221
rect 96 -549197 102 -548221
rect 56 -549209 102 -549197
rect -46 -549247 46 -549241
rect -46 -549281 -34 -549247
rect 34 -549281 46 -549247
rect -46 -549287 46 -549281
rect -46 -549355 46 -549349
rect -46 -549389 -34 -549355
rect 34 -549389 46 -549355
rect -46 -549395 46 -549389
rect -102 -549439 -56 -549427
rect -102 -550415 -96 -549439
rect -62 -550415 -56 -549439
rect -102 -550427 -56 -550415
rect 56 -549439 102 -549427
rect 56 -550415 62 -549439
rect 96 -550415 102 -549439
rect 56 -550427 102 -550415
rect -46 -550465 46 -550459
rect -46 -550499 -34 -550465
rect 34 -550499 46 -550465
rect -46 -550505 46 -550499
rect -46 -550573 46 -550567
rect -46 -550607 -34 -550573
rect 34 -550607 46 -550573
rect -46 -550613 46 -550607
rect -102 -550657 -56 -550645
rect -102 -551633 -96 -550657
rect -62 -551633 -56 -550657
rect -102 -551645 -56 -551633
rect 56 -550657 102 -550645
rect 56 -551633 62 -550657
rect 96 -551633 102 -550657
rect 56 -551645 102 -551633
rect -46 -551683 46 -551677
rect -46 -551717 -34 -551683
rect 34 -551717 46 -551683
rect -46 -551723 46 -551717
rect -46 -551791 46 -551785
rect -46 -551825 -34 -551791
rect 34 -551825 46 -551791
rect -46 -551831 46 -551825
rect -102 -551875 -56 -551863
rect -102 -552851 -96 -551875
rect -62 -552851 -56 -551875
rect -102 -552863 -56 -552851
rect 56 -551875 102 -551863
rect 56 -552851 62 -551875
rect 96 -552851 102 -551875
rect 56 -552863 102 -552851
rect -46 -552901 46 -552895
rect -46 -552935 -34 -552901
rect 34 -552935 46 -552901
rect -46 -552941 46 -552935
rect -46 -553009 46 -553003
rect -46 -553043 -34 -553009
rect 34 -553043 46 -553009
rect -46 -553049 46 -553043
rect -102 -553093 -56 -553081
rect -102 -554069 -96 -553093
rect -62 -554069 -56 -553093
rect -102 -554081 -56 -554069
rect 56 -553093 102 -553081
rect 56 -554069 62 -553093
rect 96 -554069 102 -553093
rect 56 -554081 102 -554069
rect -46 -554119 46 -554113
rect -46 -554153 -34 -554119
rect 34 -554153 46 -554119
rect -46 -554159 46 -554153
rect -46 -554227 46 -554221
rect -46 -554261 -34 -554227
rect 34 -554261 46 -554227
rect -46 -554267 46 -554261
rect -102 -554311 -56 -554299
rect -102 -555287 -96 -554311
rect -62 -555287 -56 -554311
rect -102 -555299 -56 -555287
rect 56 -554311 102 -554299
rect 56 -555287 62 -554311
rect 96 -555287 102 -554311
rect 56 -555299 102 -555287
rect -46 -555337 46 -555331
rect -46 -555371 -34 -555337
rect 34 -555371 46 -555337
rect -46 -555377 46 -555371
rect -46 -555445 46 -555439
rect -46 -555479 -34 -555445
rect 34 -555479 46 -555445
rect -46 -555485 46 -555479
rect -102 -555529 -56 -555517
rect -102 -556505 -96 -555529
rect -62 -556505 -56 -555529
rect -102 -556517 -56 -556505
rect 56 -555529 102 -555517
rect 56 -556505 62 -555529
rect 96 -556505 102 -555529
rect 56 -556517 102 -556505
rect -46 -556555 46 -556549
rect -46 -556589 -34 -556555
rect 34 -556589 46 -556555
rect -46 -556595 46 -556589
rect -46 -556663 46 -556657
rect -46 -556697 -34 -556663
rect 34 -556697 46 -556663
rect -46 -556703 46 -556697
rect -102 -556747 -56 -556735
rect -102 -557723 -96 -556747
rect -62 -557723 -56 -556747
rect -102 -557735 -56 -557723
rect 56 -556747 102 -556735
rect 56 -557723 62 -556747
rect 96 -557723 102 -556747
rect 56 -557735 102 -557723
rect -46 -557773 46 -557767
rect -46 -557807 -34 -557773
rect 34 -557807 46 -557773
rect -46 -557813 46 -557807
rect -46 -557881 46 -557875
rect -46 -557915 -34 -557881
rect 34 -557915 46 -557881
rect -46 -557921 46 -557915
rect -102 -557965 -56 -557953
rect -102 -558941 -96 -557965
rect -62 -558941 -56 -557965
rect -102 -558953 -56 -558941
rect 56 -557965 102 -557953
rect 56 -558941 62 -557965
rect 96 -558941 102 -557965
rect 56 -558953 102 -558941
rect -46 -558991 46 -558985
rect -46 -559025 -34 -558991
rect 34 -559025 46 -558991
rect -46 -559031 46 -559025
rect -46 -559099 46 -559093
rect -46 -559133 -34 -559099
rect 34 -559133 46 -559099
rect -46 -559139 46 -559133
rect -102 -559183 -56 -559171
rect -102 -560159 -96 -559183
rect -62 -560159 -56 -559183
rect -102 -560171 -56 -560159
rect 56 -559183 102 -559171
rect 56 -560159 62 -559183
rect 96 -560159 102 -559183
rect 56 -560171 102 -560159
rect -46 -560209 46 -560203
rect -46 -560243 -34 -560209
rect 34 -560243 46 -560209
rect -46 -560249 46 -560243
rect -46 -560317 46 -560311
rect -46 -560351 -34 -560317
rect 34 -560351 46 -560317
rect -46 -560357 46 -560351
rect -102 -560401 -56 -560389
rect -102 -561377 -96 -560401
rect -62 -561377 -56 -560401
rect -102 -561389 -56 -561377
rect 56 -560401 102 -560389
rect 56 -561377 62 -560401
rect 96 -561377 102 -560401
rect 56 -561389 102 -561377
rect -46 -561427 46 -561421
rect -46 -561461 -34 -561427
rect 34 -561461 46 -561427
rect -46 -561467 46 -561461
rect -46 -561535 46 -561529
rect -46 -561569 -34 -561535
rect 34 -561569 46 -561535
rect -46 -561575 46 -561569
rect -102 -561619 -56 -561607
rect -102 -562595 -96 -561619
rect -62 -562595 -56 -561619
rect -102 -562607 -56 -562595
rect 56 -561619 102 -561607
rect 56 -562595 62 -561619
rect 96 -562595 102 -561619
rect 56 -562607 102 -562595
rect -46 -562645 46 -562639
rect -46 -562679 -34 -562645
rect 34 -562679 46 -562645
rect -46 -562685 46 -562679
rect -46 -562753 46 -562747
rect -46 -562787 -34 -562753
rect 34 -562787 46 -562753
rect -46 -562793 46 -562787
rect -102 -562837 -56 -562825
rect -102 -563813 -96 -562837
rect -62 -563813 -56 -562837
rect -102 -563825 -56 -563813
rect 56 -562837 102 -562825
rect 56 -563813 62 -562837
rect 96 -563813 102 -562837
rect 56 -563825 102 -563813
rect -46 -563863 46 -563857
rect -46 -563897 -34 -563863
rect 34 -563897 46 -563863
rect -46 -563903 46 -563897
rect -46 -563971 46 -563965
rect -46 -564005 -34 -563971
rect 34 -564005 46 -563971
rect -46 -564011 46 -564005
rect -102 -564055 -56 -564043
rect -102 -565031 -96 -564055
rect -62 -565031 -56 -564055
rect -102 -565043 -56 -565031
rect 56 -564055 102 -564043
rect 56 -565031 62 -564055
rect 96 -565031 102 -564055
rect 56 -565043 102 -565031
rect -46 -565081 46 -565075
rect -46 -565115 -34 -565081
rect 34 -565115 46 -565081
rect -46 -565121 46 -565115
rect -46 -565189 46 -565183
rect -46 -565223 -34 -565189
rect 34 -565223 46 -565189
rect -46 -565229 46 -565223
rect -102 -565273 -56 -565261
rect -102 -566249 -96 -565273
rect -62 -566249 -56 -565273
rect -102 -566261 -56 -566249
rect 56 -565273 102 -565261
rect 56 -566249 62 -565273
rect 96 -566249 102 -565273
rect 56 -566261 102 -566249
rect -46 -566299 46 -566293
rect -46 -566333 -34 -566299
rect 34 -566333 46 -566299
rect -46 -566339 46 -566333
rect -46 -566407 46 -566401
rect -46 -566441 -34 -566407
rect 34 -566441 46 -566407
rect -46 -566447 46 -566441
rect -102 -566491 -56 -566479
rect -102 -567467 -96 -566491
rect -62 -567467 -56 -566491
rect -102 -567479 -56 -567467
rect 56 -566491 102 -566479
rect 56 -567467 62 -566491
rect 96 -567467 102 -566491
rect 56 -567479 102 -567467
rect -46 -567517 46 -567511
rect -46 -567551 -34 -567517
rect 34 -567551 46 -567517
rect -46 -567557 46 -567551
rect -46 -567625 46 -567619
rect -46 -567659 -34 -567625
rect 34 -567659 46 -567625
rect -46 -567665 46 -567659
rect -102 -567709 -56 -567697
rect -102 -568685 -96 -567709
rect -62 -568685 -56 -567709
rect -102 -568697 -56 -568685
rect 56 -567709 102 -567697
rect 56 -568685 62 -567709
rect 96 -568685 102 -567709
rect 56 -568697 102 -568685
rect -46 -568735 46 -568729
rect -46 -568769 -34 -568735
rect 34 -568769 46 -568735
rect -46 -568775 46 -568769
rect -46 -568843 46 -568837
rect -46 -568877 -34 -568843
rect 34 -568877 46 -568843
rect -46 -568883 46 -568877
rect -102 -568927 -56 -568915
rect -102 -569903 -96 -568927
rect -62 -569903 -56 -568927
rect -102 -569915 -56 -569903
rect 56 -568927 102 -568915
rect 56 -569903 62 -568927
rect 96 -569903 102 -568927
rect 56 -569915 102 -569903
rect -46 -569953 46 -569947
rect -46 -569987 -34 -569953
rect 34 -569987 46 -569953
rect -46 -569993 46 -569987
rect -46 -570061 46 -570055
rect -46 -570095 -34 -570061
rect 34 -570095 46 -570061
rect -46 -570101 46 -570095
rect -102 -570145 -56 -570133
rect -102 -571121 -96 -570145
rect -62 -571121 -56 -570145
rect -102 -571133 -56 -571121
rect 56 -570145 102 -570133
rect 56 -571121 62 -570145
rect 96 -571121 102 -570145
rect 56 -571133 102 -571121
rect -46 -571171 46 -571165
rect -46 -571205 -34 -571171
rect 34 -571205 46 -571171
rect -46 -571211 46 -571205
rect -46 -571279 46 -571273
rect -46 -571313 -34 -571279
rect 34 -571313 46 -571279
rect -46 -571319 46 -571313
rect -102 -571363 -56 -571351
rect -102 -572339 -96 -571363
rect -62 -572339 -56 -571363
rect -102 -572351 -56 -572339
rect 56 -571363 102 -571351
rect 56 -572339 62 -571363
rect 96 -572339 102 -571363
rect 56 -572351 102 -572339
rect -46 -572389 46 -572383
rect -46 -572423 -34 -572389
rect 34 -572423 46 -572389
rect -46 -572429 46 -572423
rect -46 -572497 46 -572491
rect -46 -572531 -34 -572497
rect 34 -572531 46 -572497
rect -46 -572537 46 -572531
rect -102 -572581 -56 -572569
rect -102 -573557 -96 -572581
rect -62 -573557 -56 -572581
rect -102 -573569 -56 -573557
rect 56 -572581 102 -572569
rect 56 -573557 62 -572581
rect 96 -573557 102 -572581
rect 56 -573569 102 -573557
rect -46 -573607 46 -573601
rect -46 -573641 -34 -573607
rect 34 -573641 46 -573607
rect -46 -573647 46 -573641
rect -46 -573715 46 -573709
rect -46 -573749 -34 -573715
rect 34 -573749 46 -573715
rect -46 -573755 46 -573749
rect -102 -573799 -56 -573787
rect -102 -574775 -96 -573799
rect -62 -574775 -56 -573799
rect -102 -574787 -56 -574775
rect 56 -573799 102 -573787
rect 56 -574775 62 -573799
rect 96 -574775 102 -573799
rect 56 -574787 102 -574775
rect -46 -574825 46 -574819
rect -46 -574859 -34 -574825
rect 34 -574859 46 -574825
rect -46 -574865 46 -574859
rect -46 -574933 46 -574927
rect -46 -574967 -34 -574933
rect 34 -574967 46 -574933
rect -46 -574973 46 -574967
rect -102 -575017 -56 -575005
rect -102 -575993 -96 -575017
rect -62 -575993 -56 -575017
rect -102 -576005 -56 -575993
rect 56 -575017 102 -575005
rect 56 -575993 62 -575017
rect 96 -575993 102 -575017
rect 56 -576005 102 -575993
rect -46 -576043 46 -576037
rect -46 -576077 -34 -576043
rect 34 -576077 46 -576043
rect -46 -576083 46 -576077
rect -46 -576151 46 -576145
rect -46 -576185 -34 -576151
rect 34 -576185 46 -576151
rect -46 -576191 46 -576185
rect -102 -576235 -56 -576223
rect -102 -577211 -96 -576235
rect -62 -577211 -56 -576235
rect -102 -577223 -56 -577211
rect 56 -576235 102 -576223
rect 56 -577211 62 -576235
rect 96 -577211 102 -576235
rect 56 -577223 102 -577211
rect -46 -577261 46 -577255
rect -46 -577295 -34 -577261
rect 34 -577295 46 -577261
rect -46 -577301 46 -577295
rect -46 -577369 46 -577363
rect -46 -577403 -34 -577369
rect 34 -577403 46 -577369
rect -46 -577409 46 -577403
rect -102 -577453 -56 -577441
rect -102 -578429 -96 -577453
rect -62 -578429 -56 -577453
rect -102 -578441 -56 -578429
rect 56 -577453 102 -577441
rect 56 -578429 62 -577453
rect 96 -578429 102 -577453
rect 56 -578441 102 -578429
rect -46 -578479 46 -578473
rect -46 -578513 -34 -578479
rect 34 -578513 46 -578479
rect -46 -578519 46 -578513
rect -46 -578587 46 -578581
rect -46 -578621 -34 -578587
rect 34 -578621 46 -578587
rect -46 -578627 46 -578621
rect -102 -578671 -56 -578659
rect -102 -579647 -96 -578671
rect -62 -579647 -56 -578671
rect -102 -579659 -56 -579647
rect 56 -578671 102 -578659
rect 56 -579647 62 -578671
rect 96 -579647 102 -578671
rect 56 -579659 102 -579647
rect -46 -579697 46 -579691
rect -46 -579731 -34 -579697
rect 34 -579731 46 -579697
rect -46 -579737 46 -579731
rect -46 -579805 46 -579799
rect -46 -579839 -34 -579805
rect 34 -579839 46 -579805
rect -46 -579845 46 -579839
rect -102 -579889 -56 -579877
rect -102 -580865 -96 -579889
rect -62 -580865 -56 -579889
rect -102 -580877 -56 -580865
rect 56 -579889 102 -579877
rect 56 -580865 62 -579889
rect 96 -580865 102 -579889
rect 56 -580877 102 -580865
rect -46 -580915 46 -580909
rect -46 -580949 -34 -580915
rect 34 -580949 46 -580915
rect -46 -580955 46 -580949
rect -46 -581023 46 -581017
rect -46 -581057 -34 -581023
rect 34 -581057 46 -581023
rect -46 -581063 46 -581057
rect -102 -581107 -56 -581095
rect -102 -582083 -96 -581107
rect -62 -582083 -56 -581107
rect -102 -582095 -56 -582083
rect 56 -581107 102 -581095
rect 56 -582083 62 -581107
rect 96 -582083 102 -581107
rect 56 -582095 102 -582083
rect -46 -582133 46 -582127
rect -46 -582167 -34 -582133
rect 34 -582167 46 -582133
rect -46 -582173 46 -582167
rect -46 -582241 46 -582235
rect -46 -582275 -34 -582241
rect 34 -582275 46 -582241
rect -46 -582281 46 -582275
rect -102 -582325 -56 -582313
rect -102 -583301 -96 -582325
rect -62 -583301 -56 -582325
rect -102 -583313 -56 -583301
rect 56 -582325 102 -582313
rect 56 -583301 62 -582325
rect 96 -583301 102 -582325
rect 56 -583313 102 -583301
rect -46 -583351 46 -583345
rect -46 -583385 -34 -583351
rect 34 -583385 46 -583351
rect -46 -583391 46 -583385
rect -46 -583459 46 -583453
rect -46 -583493 -34 -583459
rect 34 -583493 46 -583459
rect -46 -583499 46 -583493
rect -102 -583543 -56 -583531
rect -102 -584519 -96 -583543
rect -62 -584519 -56 -583543
rect -102 -584531 -56 -584519
rect 56 -583543 102 -583531
rect 56 -584519 62 -583543
rect 96 -584519 102 -583543
rect 56 -584531 102 -584519
rect -46 -584569 46 -584563
rect -46 -584603 -34 -584569
rect 34 -584603 46 -584569
rect -46 -584609 46 -584603
rect -46 -584677 46 -584671
rect -46 -584711 -34 -584677
rect 34 -584711 46 -584677
rect -46 -584717 46 -584711
rect -102 -584761 -56 -584749
rect -102 -585737 -96 -584761
rect -62 -585737 -56 -584761
rect -102 -585749 -56 -585737
rect 56 -584761 102 -584749
rect 56 -585737 62 -584761
rect 96 -585737 102 -584761
rect 56 -585749 102 -585737
rect -46 -585787 46 -585781
rect -46 -585821 -34 -585787
rect 34 -585821 46 -585787
rect -46 -585827 46 -585821
rect -46 -585895 46 -585889
rect -46 -585929 -34 -585895
rect 34 -585929 46 -585895
rect -46 -585935 46 -585929
rect -102 -585979 -56 -585967
rect -102 -586955 -96 -585979
rect -62 -586955 -56 -585979
rect -102 -586967 -56 -586955
rect 56 -585979 102 -585967
rect 56 -586955 62 -585979
rect 96 -586955 102 -585979
rect 56 -586967 102 -586955
rect -46 -587005 46 -586999
rect -46 -587039 -34 -587005
rect 34 -587039 46 -587005
rect -46 -587045 46 -587039
rect -46 -587113 46 -587107
rect -46 -587147 -34 -587113
rect 34 -587147 46 -587113
rect -46 -587153 46 -587147
rect -102 -587197 -56 -587185
rect -102 -588173 -96 -587197
rect -62 -588173 -56 -587197
rect -102 -588185 -56 -588173
rect 56 -587197 102 -587185
rect 56 -588173 62 -587197
rect 96 -588173 102 -587197
rect 56 -588185 102 -588173
rect -46 -588223 46 -588217
rect -46 -588257 -34 -588223
rect 34 -588257 46 -588223
rect -46 -588263 46 -588257
rect -46 -588331 46 -588325
rect -46 -588365 -34 -588331
rect 34 -588365 46 -588331
rect -46 -588371 46 -588365
rect -102 -588415 -56 -588403
rect -102 -589391 -96 -588415
rect -62 -589391 -56 -588415
rect -102 -589403 -56 -589391
rect 56 -588415 102 -588403
rect 56 -589391 62 -588415
rect 96 -589391 102 -588415
rect 56 -589403 102 -589391
rect -46 -589441 46 -589435
rect -46 -589475 -34 -589441
rect 34 -589475 46 -589441
rect -46 -589481 46 -589475
rect -46 -589549 46 -589543
rect -46 -589583 -34 -589549
rect 34 -589583 46 -589549
rect -46 -589589 46 -589583
rect -102 -589633 -56 -589621
rect -102 -590609 -96 -589633
rect -62 -590609 -56 -589633
rect -102 -590621 -56 -590609
rect 56 -589633 102 -589621
rect 56 -590609 62 -589633
rect 96 -590609 102 -589633
rect 56 -590621 102 -590609
rect -46 -590659 46 -590653
rect -46 -590693 -34 -590659
rect 34 -590693 46 -590659
rect -46 -590699 46 -590693
rect -46 -590767 46 -590761
rect -46 -590801 -34 -590767
rect 34 -590801 46 -590767
rect -46 -590807 46 -590801
rect -102 -590851 -56 -590839
rect -102 -591827 -96 -590851
rect -62 -591827 -56 -590851
rect -102 -591839 -56 -591827
rect 56 -590851 102 -590839
rect 56 -591827 62 -590851
rect 96 -591827 102 -590851
rect 56 -591839 102 -591827
rect -46 -591877 46 -591871
rect -46 -591911 -34 -591877
rect 34 -591911 46 -591877
rect -46 -591917 46 -591911
rect -46 -591985 46 -591979
rect -46 -592019 -34 -591985
rect 34 -592019 46 -591985
rect -46 -592025 46 -592019
rect -102 -592069 -56 -592057
rect -102 -593045 -96 -592069
rect -62 -593045 -56 -592069
rect -102 -593057 -56 -593045
rect 56 -592069 102 -592057
rect 56 -593045 62 -592069
rect 96 -593045 102 -592069
rect 56 -593057 102 -593045
rect -46 -593095 46 -593089
rect -46 -593129 -34 -593095
rect 34 -593129 46 -593095
rect -46 -593135 46 -593129
rect -46 -593203 46 -593197
rect -46 -593237 -34 -593203
rect 34 -593237 46 -593203
rect -46 -593243 46 -593237
rect -102 -593287 -56 -593275
rect -102 -594263 -96 -593287
rect -62 -594263 -56 -593287
rect -102 -594275 -56 -594263
rect 56 -593287 102 -593275
rect 56 -594263 62 -593287
rect 96 -594263 102 -593287
rect 56 -594275 102 -594263
rect -46 -594313 46 -594307
rect -46 -594347 -34 -594313
rect 34 -594347 46 -594313
rect -46 -594353 46 -594347
rect -46 -594421 46 -594415
rect -46 -594455 -34 -594421
rect 34 -594455 46 -594421
rect -46 -594461 46 -594455
rect -102 -594505 -56 -594493
rect -102 -595481 -96 -594505
rect -62 -595481 -56 -594505
rect -102 -595493 -56 -595481
rect 56 -594505 102 -594493
rect 56 -595481 62 -594505
rect 96 -595481 102 -594505
rect 56 -595493 102 -595481
rect -46 -595531 46 -595525
rect -46 -595565 -34 -595531
rect 34 -595565 46 -595531
rect -46 -595571 46 -595565
rect -46 -595639 46 -595633
rect -46 -595673 -34 -595639
rect 34 -595673 46 -595639
rect -46 -595679 46 -595673
rect -102 -595723 -56 -595711
rect -102 -596699 -96 -595723
rect -62 -596699 -56 -595723
rect -102 -596711 -56 -596699
rect 56 -595723 102 -595711
rect 56 -596699 62 -595723
rect 96 -596699 102 -595723
rect 56 -596711 102 -596699
rect -46 -596749 46 -596743
rect -46 -596783 -34 -596749
rect 34 -596783 46 -596749
rect -46 -596789 46 -596783
rect -46 -596857 46 -596851
rect -46 -596891 -34 -596857
rect 34 -596891 46 -596857
rect -46 -596897 46 -596891
rect -102 -596941 -56 -596929
rect -102 -597917 -96 -596941
rect -62 -597917 -56 -596941
rect -102 -597929 -56 -597917
rect 56 -596941 102 -596929
rect 56 -597917 62 -596941
rect 96 -597917 102 -596941
rect 56 -597929 102 -597917
rect -46 -597967 46 -597961
rect -46 -598001 -34 -597967
rect 34 -598001 46 -597967
rect -46 -598007 46 -598001
rect -46 -598075 46 -598069
rect -46 -598109 -34 -598075
rect 34 -598109 46 -598075
rect -46 -598115 46 -598109
rect -102 -598159 -56 -598147
rect -102 -599135 -96 -598159
rect -62 -599135 -56 -598159
rect -102 -599147 -56 -599135
rect 56 -598159 102 -598147
rect 56 -599135 62 -598159
rect 96 -599135 102 -598159
rect 56 -599147 102 -599135
rect -46 -599185 46 -599179
rect -46 -599219 -34 -599185
rect 34 -599219 46 -599185
rect -46 -599225 46 -599219
rect -46 -599293 46 -599287
rect -46 -599327 -34 -599293
rect 34 -599327 46 -599293
rect -46 -599333 46 -599327
rect -102 -599377 -56 -599365
rect -102 -600353 -96 -599377
rect -62 -600353 -56 -599377
rect -102 -600365 -56 -600353
rect 56 -599377 102 -599365
rect 56 -600353 62 -599377
rect 96 -600353 102 -599377
rect 56 -600365 102 -600353
rect -46 -600403 46 -600397
rect -46 -600437 -34 -600403
rect 34 -600437 46 -600403
rect -46 -600443 46 -600437
rect -46 -600511 46 -600505
rect -46 -600545 -34 -600511
rect 34 -600545 46 -600511
rect -46 -600551 46 -600545
rect -102 -600595 -56 -600583
rect -102 -601571 -96 -600595
rect -62 -601571 -56 -600595
rect -102 -601583 -56 -601571
rect 56 -600595 102 -600583
rect 56 -601571 62 -600595
rect 96 -601571 102 -600595
rect 56 -601583 102 -601571
rect -46 -601621 46 -601615
rect -46 -601655 -34 -601621
rect 34 -601655 46 -601621
rect -46 -601661 46 -601655
rect -46 -601729 46 -601723
rect -46 -601763 -34 -601729
rect 34 -601763 46 -601729
rect -46 -601769 46 -601763
rect -102 -601813 -56 -601801
rect -102 -602789 -96 -601813
rect -62 -602789 -56 -601813
rect -102 -602801 -56 -602789
rect 56 -601813 102 -601801
rect 56 -602789 62 -601813
rect 96 -602789 102 -601813
rect 56 -602801 102 -602789
rect -46 -602839 46 -602833
rect -46 -602873 -34 -602839
rect 34 -602873 46 -602839
rect -46 -602879 46 -602873
rect -46 -602947 46 -602941
rect -46 -602981 -34 -602947
rect 34 -602981 46 -602947
rect -46 -602987 46 -602981
rect -102 -603031 -56 -603019
rect -102 -604007 -96 -603031
rect -62 -604007 -56 -603031
rect -102 -604019 -56 -604007
rect 56 -603031 102 -603019
rect 56 -604007 62 -603031
rect 96 -604007 102 -603031
rect 56 -604019 102 -604007
rect -46 -604057 46 -604051
rect -46 -604091 -34 -604057
rect 34 -604091 46 -604057
rect -46 -604097 46 -604091
rect -46 -604165 46 -604159
rect -46 -604199 -34 -604165
rect 34 -604199 46 -604165
rect -46 -604205 46 -604199
rect -102 -604249 -56 -604237
rect -102 -605225 -96 -604249
rect -62 -605225 -56 -604249
rect -102 -605237 -56 -605225
rect 56 -604249 102 -604237
rect 56 -605225 62 -604249
rect 96 -605225 102 -604249
rect 56 -605237 102 -605225
rect -46 -605275 46 -605269
rect -46 -605309 -34 -605275
rect 34 -605309 46 -605275
rect -46 -605315 46 -605309
rect -46 -605383 46 -605377
rect -46 -605417 -34 -605383
rect 34 -605417 46 -605383
rect -46 -605423 46 -605417
rect -102 -605467 -56 -605455
rect -102 -606443 -96 -605467
rect -62 -606443 -56 -605467
rect -102 -606455 -56 -606443
rect 56 -605467 102 -605455
rect 56 -606443 62 -605467
rect 96 -606443 102 -605467
rect 56 -606455 102 -606443
rect -46 -606493 46 -606487
rect -46 -606527 -34 -606493
rect 34 -606527 46 -606493
rect -46 -606533 46 -606527
rect -46 -606601 46 -606595
rect -46 -606635 -34 -606601
rect 34 -606635 46 -606601
rect -46 -606641 46 -606635
rect -102 -606685 -56 -606673
rect -102 -607661 -96 -606685
rect -62 -607661 -56 -606685
rect -102 -607673 -56 -607661
rect 56 -606685 102 -606673
rect 56 -607661 62 -606685
rect 96 -607661 102 -606685
rect 56 -607673 102 -607661
rect -46 -607711 46 -607705
rect -46 -607745 -34 -607711
rect 34 -607745 46 -607711
rect -46 -607751 46 -607745
rect -46 -607819 46 -607813
rect -46 -607853 -34 -607819
rect 34 -607853 46 -607819
rect -46 -607859 46 -607853
rect -102 -607903 -56 -607891
rect -102 -608879 -96 -607903
rect -62 -608879 -56 -607903
rect -102 -608891 -56 -608879
rect 56 -607903 102 -607891
rect 56 -608879 62 -607903
rect 96 -608879 102 -607903
rect 56 -608891 102 -608879
rect -46 -608929 46 -608923
rect -46 -608963 -34 -608929
rect 34 -608963 46 -608929
rect -46 -608969 46 -608963
<< properties >>
string FIXED_BBOX -213 -609084 213 609084
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1000 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
