magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< nwell >>
rect -1258 -1269 1258 1269
<< mvpmos >>
rect -1000 772 1000 972
rect -1000 336 1000 536
rect -1000 -100 1000 100
rect -1000 -536 1000 -336
rect -1000 -972 1000 -772
<< mvpdiff >>
rect -1058 960 -1000 972
rect -1058 784 -1046 960
rect -1012 784 -1000 960
rect -1058 772 -1000 784
rect 1000 960 1058 972
rect 1000 784 1012 960
rect 1046 784 1058 960
rect 1000 772 1058 784
rect -1058 524 -1000 536
rect -1058 348 -1046 524
rect -1012 348 -1000 524
rect -1058 336 -1000 348
rect 1000 524 1058 536
rect 1000 348 1012 524
rect 1046 348 1058 524
rect 1000 336 1058 348
rect -1058 88 -1000 100
rect -1058 -88 -1046 88
rect -1012 -88 -1000 88
rect -1058 -100 -1000 -88
rect 1000 88 1058 100
rect 1000 -88 1012 88
rect 1046 -88 1058 88
rect 1000 -100 1058 -88
rect -1058 -348 -1000 -336
rect -1058 -524 -1046 -348
rect -1012 -524 -1000 -348
rect -1058 -536 -1000 -524
rect 1000 -348 1058 -336
rect 1000 -524 1012 -348
rect 1046 -524 1058 -348
rect 1000 -536 1058 -524
rect -1058 -784 -1000 -772
rect -1058 -960 -1046 -784
rect -1012 -960 -1000 -784
rect -1058 -972 -1000 -960
rect 1000 -784 1058 -772
rect 1000 -960 1012 -784
rect 1046 -960 1058 -784
rect 1000 -972 1058 -960
<< mvpdiffc >>
rect -1046 784 -1012 960
rect 1012 784 1046 960
rect -1046 348 -1012 524
rect 1012 348 1046 524
rect -1046 -88 -1012 88
rect 1012 -88 1046 88
rect -1046 -524 -1012 -348
rect 1012 -524 1046 -348
rect -1046 -960 -1012 -784
rect 1012 -960 1046 -784
<< mvnsubdiff >>
rect -1192 1191 1192 1203
rect -1192 1157 -1084 1191
rect 1084 1157 1192 1191
rect -1192 1145 1192 1157
rect -1192 1095 -1134 1145
rect -1192 -1095 -1180 1095
rect -1146 -1095 -1134 1095
rect 1134 1095 1192 1145
rect -1192 -1145 -1134 -1095
rect 1134 -1095 1146 1095
rect 1180 -1095 1192 1095
rect 1134 -1145 1192 -1095
rect -1192 -1157 1192 -1145
rect -1192 -1191 -1084 -1157
rect 1084 -1191 1192 -1157
rect -1192 -1203 1192 -1191
<< mvnsubdiffcont >>
rect -1084 1157 1084 1191
rect -1180 -1095 -1146 1095
rect 1146 -1095 1180 1095
rect -1084 -1191 1084 -1157
<< poly >>
rect -1000 1053 1000 1069
rect -1000 1019 -984 1053
rect 984 1019 1000 1053
rect -1000 972 1000 1019
rect -1000 725 1000 772
rect -1000 691 -984 725
rect 984 691 1000 725
rect -1000 675 1000 691
rect -1000 617 1000 633
rect -1000 583 -984 617
rect 984 583 1000 617
rect -1000 536 1000 583
rect -1000 289 1000 336
rect -1000 255 -984 289
rect 984 255 1000 289
rect -1000 239 1000 255
rect -1000 181 1000 197
rect -1000 147 -984 181
rect 984 147 1000 181
rect -1000 100 1000 147
rect -1000 -147 1000 -100
rect -1000 -181 -984 -147
rect 984 -181 1000 -147
rect -1000 -197 1000 -181
rect -1000 -255 1000 -239
rect -1000 -289 -984 -255
rect 984 -289 1000 -255
rect -1000 -336 1000 -289
rect -1000 -583 1000 -536
rect -1000 -617 -984 -583
rect 984 -617 1000 -583
rect -1000 -633 1000 -617
rect -1000 -691 1000 -675
rect -1000 -725 -984 -691
rect 984 -725 1000 -691
rect -1000 -772 1000 -725
rect -1000 -1019 1000 -972
rect -1000 -1053 -984 -1019
rect 984 -1053 1000 -1019
rect -1000 -1069 1000 -1053
<< polycont >>
rect -984 1019 984 1053
rect -984 691 984 725
rect -984 583 984 617
rect -984 255 984 289
rect -984 147 984 181
rect -984 -181 984 -147
rect -984 -289 984 -255
rect -984 -617 984 -583
rect -984 -725 984 -691
rect -984 -1053 984 -1019
<< locali >>
rect -1180 1157 -1084 1191
rect 1084 1157 1180 1191
rect -1180 1095 -1146 1157
rect 1146 1095 1180 1157
rect -1000 1019 -984 1053
rect 984 1019 1000 1053
rect -1046 960 -1012 976
rect -1046 768 -1012 784
rect 1012 960 1046 976
rect 1012 768 1046 784
rect -1000 691 -984 725
rect 984 691 1000 725
rect -1000 583 -984 617
rect 984 583 1000 617
rect -1046 524 -1012 540
rect -1046 332 -1012 348
rect 1012 524 1046 540
rect 1012 332 1046 348
rect -1000 255 -984 289
rect 984 255 1000 289
rect -1000 147 -984 181
rect 984 147 1000 181
rect -1046 88 -1012 104
rect -1046 -104 -1012 -88
rect 1012 88 1046 104
rect 1012 -104 1046 -88
rect -1000 -181 -984 -147
rect 984 -181 1000 -147
rect -1000 -289 -984 -255
rect 984 -289 1000 -255
rect -1046 -348 -1012 -332
rect -1046 -540 -1012 -524
rect 1012 -348 1046 -332
rect 1012 -540 1046 -524
rect -1000 -617 -984 -583
rect 984 -617 1000 -583
rect -1000 -725 -984 -691
rect 984 -725 1000 -691
rect -1046 -784 -1012 -768
rect -1046 -976 -1012 -960
rect 1012 -784 1046 -768
rect 1012 -976 1046 -960
rect -1000 -1053 -984 -1019
rect 984 -1053 1000 -1019
rect -1180 -1157 -1146 -1095
rect 1146 -1157 1180 -1095
rect -1180 -1191 -1084 -1157
rect 1084 -1191 1180 -1157
<< viali >>
rect -984 1019 984 1053
rect -1046 784 -1012 960
rect 1012 784 1046 960
rect -984 691 984 725
rect -984 583 984 617
rect -1046 348 -1012 524
rect 1012 348 1046 524
rect -984 255 984 289
rect -984 147 984 181
rect -1046 -88 -1012 88
rect 1012 -88 1046 88
rect -984 -181 984 -147
rect -984 -289 984 -255
rect -1046 -524 -1012 -348
rect 1012 -524 1046 -348
rect -984 -617 984 -583
rect -984 -725 984 -691
rect -1046 -960 -1012 -784
rect 1012 -960 1046 -784
rect -984 -1053 984 -1019
<< metal1 >>
rect -996 1053 996 1059
rect -996 1019 -984 1053
rect 984 1019 996 1053
rect -996 1013 996 1019
rect -1052 960 -1006 972
rect -1052 784 -1046 960
rect -1012 784 -1006 960
rect -1052 772 -1006 784
rect 1006 960 1052 972
rect 1006 784 1012 960
rect 1046 784 1052 960
rect 1006 772 1052 784
rect -996 725 996 731
rect -996 691 -984 725
rect 984 691 996 725
rect -996 685 996 691
rect -996 617 996 623
rect -996 583 -984 617
rect 984 583 996 617
rect -996 577 996 583
rect -1052 524 -1006 536
rect -1052 348 -1046 524
rect -1012 348 -1006 524
rect -1052 336 -1006 348
rect 1006 524 1052 536
rect 1006 348 1012 524
rect 1046 348 1052 524
rect 1006 336 1052 348
rect -996 289 996 295
rect -996 255 -984 289
rect 984 255 996 289
rect -996 249 996 255
rect -996 181 996 187
rect -996 147 -984 181
rect 984 147 996 181
rect -996 141 996 147
rect -1052 88 -1006 100
rect -1052 -88 -1046 88
rect -1012 -88 -1006 88
rect -1052 -100 -1006 -88
rect 1006 88 1052 100
rect 1006 -88 1012 88
rect 1046 -88 1052 88
rect 1006 -100 1052 -88
rect -996 -147 996 -141
rect -996 -181 -984 -147
rect 984 -181 996 -147
rect -996 -187 996 -181
rect -996 -255 996 -249
rect -996 -289 -984 -255
rect 984 -289 996 -255
rect -996 -295 996 -289
rect -1052 -348 -1006 -336
rect -1052 -524 -1046 -348
rect -1012 -524 -1006 -348
rect -1052 -536 -1006 -524
rect 1006 -348 1052 -336
rect 1006 -524 1012 -348
rect 1046 -524 1052 -348
rect 1006 -536 1052 -524
rect -996 -583 996 -577
rect -996 -617 -984 -583
rect 984 -617 996 -583
rect -996 -623 996 -617
rect -996 -691 996 -685
rect -996 -725 -984 -691
rect 984 -725 996 -691
rect -996 -731 996 -725
rect -1052 -784 -1006 -772
rect -1052 -960 -1046 -784
rect -1012 -960 -1006 -784
rect -1052 -972 -1006 -960
rect 1006 -784 1052 -772
rect 1006 -960 1012 -784
rect 1046 -960 1052 -784
rect 1006 -972 1052 -960
rect -996 -1019 996 -1013
rect -996 -1053 -984 -1019
rect 984 -1053 996 -1019
rect -996 -1059 996 -1053
<< properties >>
string FIXED_BBOX -1163 -1174 1163 1174
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
