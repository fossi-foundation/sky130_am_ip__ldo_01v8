magic
tech sky130A
timestamp 1717294357
<< pwell >>
rect -569 -597 569 597
<< mvnmos >>
rect -450 368 450 468
rect -450 159 450 259
rect -450 -50 450 50
rect -450 -259 450 -159
rect -450 -468 450 -368
<< mvndiff >>
rect -479 462 -450 468
rect -479 374 -473 462
rect -456 374 -450 462
rect -479 368 -450 374
rect 450 462 479 468
rect 450 374 456 462
rect 473 374 479 462
rect 450 368 479 374
rect -479 253 -450 259
rect -479 165 -473 253
rect -456 165 -450 253
rect -479 159 -450 165
rect 450 253 479 259
rect 450 165 456 253
rect 473 165 479 253
rect 450 159 479 165
rect -479 44 -450 50
rect -479 -44 -473 44
rect -456 -44 -450 44
rect -479 -50 -450 -44
rect 450 44 479 50
rect 450 -44 456 44
rect 473 -44 479 44
rect 450 -50 479 -44
rect -479 -165 -450 -159
rect -479 -253 -473 -165
rect -456 -253 -450 -165
rect -479 -259 -450 -253
rect 450 -165 479 -159
rect 450 -253 456 -165
rect 473 -253 479 -165
rect 450 -259 479 -253
rect -479 -374 -450 -368
rect -479 -462 -473 -374
rect -456 -462 -450 -374
rect -479 -468 -450 -462
rect 450 -374 479 -368
rect 450 -462 456 -374
rect 473 -462 479 -374
rect 450 -468 479 -462
<< mvndiffc >>
rect -473 374 -456 462
rect 456 374 473 462
rect -473 165 -456 253
rect 456 165 473 253
rect -473 -44 -456 44
rect 456 -44 473 44
rect -473 -253 -456 -165
rect 456 -253 473 -165
rect -473 -462 -456 -374
rect 456 -462 473 -374
<< mvpsubdiff >>
rect -551 573 551 579
rect -551 556 -497 573
rect 497 556 551 573
rect -551 550 551 556
rect -551 525 -522 550
rect -551 -525 -545 525
rect -528 -525 -522 525
rect 522 525 551 550
rect -551 -550 -522 -525
rect 522 -525 528 525
rect 545 -525 551 525
rect 522 -550 551 -525
rect -551 -556 551 -550
rect -551 -573 -497 -556
rect 497 -573 551 -556
rect -551 -579 551 -573
<< mvpsubdiffcont >>
rect -497 556 497 573
rect -545 -525 -528 525
rect 528 -525 545 525
rect -497 -573 497 -556
<< poly >>
rect -450 504 450 512
rect -450 487 -442 504
rect 442 487 450 504
rect -450 468 450 487
rect -450 349 450 368
rect -450 332 -442 349
rect 442 332 450 349
rect -450 324 450 332
rect -450 295 450 303
rect -450 278 -442 295
rect 442 278 450 295
rect -450 259 450 278
rect -450 140 450 159
rect -450 123 -442 140
rect 442 123 450 140
rect -450 115 450 123
rect -450 86 450 94
rect -450 69 -442 86
rect 442 69 450 86
rect -450 50 450 69
rect -450 -69 450 -50
rect -450 -86 -442 -69
rect 442 -86 450 -69
rect -450 -94 450 -86
rect -450 -123 450 -115
rect -450 -140 -442 -123
rect 442 -140 450 -123
rect -450 -159 450 -140
rect -450 -278 450 -259
rect -450 -295 -442 -278
rect 442 -295 450 -278
rect -450 -303 450 -295
rect -450 -332 450 -324
rect -450 -349 -442 -332
rect 442 -349 450 -332
rect -450 -368 450 -349
rect -450 -487 450 -468
rect -450 -504 -442 -487
rect 442 -504 450 -487
rect -450 -512 450 -504
<< polycont >>
rect -442 487 442 504
rect -442 332 442 349
rect -442 278 442 295
rect -442 123 442 140
rect -442 69 442 86
rect -442 -86 442 -69
rect -442 -140 442 -123
rect -442 -295 442 -278
rect -442 -349 442 -332
rect -442 -504 442 -487
<< locali >>
rect -545 556 -497 573
rect 497 556 545 573
rect -545 525 -528 556
rect 528 525 545 556
rect -450 487 -442 504
rect 442 487 450 504
rect -473 462 -456 470
rect -473 366 -456 374
rect 456 462 473 470
rect 456 366 473 374
rect -450 332 -442 349
rect 442 332 450 349
rect -450 278 -442 295
rect 442 278 450 295
rect -473 253 -456 261
rect -473 157 -456 165
rect 456 253 473 261
rect 456 157 473 165
rect -450 123 -442 140
rect 442 123 450 140
rect -450 69 -442 86
rect 442 69 450 86
rect -473 44 -456 52
rect -473 -52 -456 -44
rect 456 44 473 52
rect 456 -52 473 -44
rect -450 -86 -442 -69
rect 442 -86 450 -69
rect -450 -140 -442 -123
rect 442 -140 450 -123
rect -473 -165 -456 -157
rect -473 -261 -456 -253
rect 456 -165 473 -157
rect 456 -261 473 -253
rect -450 -295 -442 -278
rect 442 -295 450 -278
rect -450 -349 -442 -332
rect 442 -349 450 -332
rect -473 -374 -456 -366
rect -473 -470 -456 -462
rect 456 -374 473 -366
rect 456 -470 473 -462
rect -450 -504 -442 -487
rect 442 -504 450 -487
rect -545 -556 -528 -525
rect 528 -556 545 -525
rect -545 -573 -497 -556
rect 497 -573 545 -556
<< viali >>
rect -442 487 442 504
rect -473 374 -456 462
rect 456 374 473 462
rect -442 332 442 349
rect -442 278 442 295
rect -473 165 -456 253
rect 456 165 473 253
rect -442 123 442 140
rect -442 69 442 86
rect -473 -44 -456 44
rect 456 -44 473 44
rect -442 -86 442 -69
rect -442 -140 442 -123
rect -473 -253 -456 -165
rect 456 -253 473 -165
rect -442 -295 442 -278
rect -442 -349 442 -332
rect -473 -462 -456 -374
rect 456 -462 473 -374
rect -442 -504 442 -487
<< metal1 >>
rect -448 504 448 507
rect -448 487 -442 504
rect 442 487 448 504
rect -448 484 448 487
rect -476 462 -453 468
rect -476 374 -473 462
rect -456 374 -453 462
rect -476 368 -453 374
rect 453 462 476 468
rect 453 374 456 462
rect 473 374 476 462
rect 453 368 476 374
rect -448 349 448 352
rect -448 332 -442 349
rect 442 332 448 349
rect -448 329 448 332
rect -448 295 448 298
rect -448 278 -442 295
rect 442 278 448 295
rect -448 275 448 278
rect -476 253 -453 259
rect -476 165 -473 253
rect -456 165 -453 253
rect -476 159 -453 165
rect 453 253 476 259
rect 453 165 456 253
rect 473 165 476 253
rect 453 159 476 165
rect -448 140 448 143
rect -448 123 -442 140
rect 442 123 448 140
rect -448 120 448 123
rect -448 86 448 89
rect -448 69 -442 86
rect 442 69 448 86
rect -448 66 448 69
rect -476 44 -453 50
rect -476 -44 -473 44
rect -456 -44 -453 44
rect -476 -50 -453 -44
rect 453 44 476 50
rect 453 -44 456 44
rect 473 -44 476 44
rect 453 -50 476 -44
rect -448 -69 448 -66
rect -448 -86 -442 -69
rect 442 -86 448 -69
rect -448 -89 448 -86
rect -448 -123 448 -120
rect -448 -140 -442 -123
rect 442 -140 448 -123
rect -448 -143 448 -140
rect -476 -165 -453 -159
rect -476 -253 -473 -165
rect -456 -253 -453 -165
rect -476 -259 -453 -253
rect 453 -165 476 -159
rect 453 -253 456 -165
rect 473 -253 476 -165
rect 453 -259 476 -253
rect -448 -278 448 -275
rect -448 -295 -442 -278
rect 442 -295 448 -278
rect -448 -298 448 -295
rect -448 -332 448 -329
rect -448 -349 -442 -332
rect 442 -349 448 -332
rect -448 -352 448 -349
rect -476 -374 -453 -368
rect -476 -462 -473 -374
rect -456 -462 -453 -374
rect -476 -468 -453 -462
rect 453 -374 476 -368
rect 453 -462 456 -374
rect 473 -462 476 -374
rect 453 -468 476 -462
rect -448 -487 448 -484
rect -448 -504 -442 -487
rect 442 -504 448 -487
rect -448 -507 448 -504
<< properties >>
string FIXED_BBOX -531 -564 531 564
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 9.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
