magic
tech sky130A
magscale 1 2
timestamp 1713186496
<< pwell >>
rect -1228 -985 1228 985
<< mvnmos >>
rect -1000 527 1000 727
rect -1000 109 1000 309
rect -1000 -309 1000 -109
rect -1000 -727 1000 -527
<< mvndiff >>
rect -1058 715 -1000 727
rect -1058 539 -1046 715
rect -1012 539 -1000 715
rect -1058 527 -1000 539
rect 1000 715 1058 727
rect 1000 539 1012 715
rect 1046 539 1058 715
rect 1000 527 1058 539
rect -1058 297 -1000 309
rect -1058 121 -1046 297
rect -1012 121 -1000 297
rect -1058 109 -1000 121
rect 1000 297 1058 309
rect 1000 121 1012 297
rect 1046 121 1058 297
rect 1000 109 1058 121
rect -1058 -121 -1000 -109
rect -1058 -297 -1046 -121
rect -1012 -297 -1000 -121
rect -1058 -309 -1000 -297
rect 1000 -121 1058 -109
rect 1000 -297 1012 -121
rect 1046 -297 1058 -121
rect 1000 -309 1058 -297
rect -1058 -539 -1000 -527
rect -1058 -715 -1046 -539
rect -1012 -715 -1000 -539
rect -1058 -727 -1000 -715
rect 1000 -539 1058 -527
rect 1000 -715 1012 -539
rect 1046 -715 1058 -539
rect 1000 -727 1058 -715
<< mvndiffc >>
rect -1046 539 -1012 715
rect 1012 539 1046 715
rect -1046 121 -1012 297
rect 1012 121 1046 297
rect -1046 -297 -1012 -121
rect 1012 -297 1046 -121
rect -1046 -715 -1012 -539
rect 1012 -715 1046 -539
<< mvpsubdiff >>
rect -1192 937 1192 949
rect -1192 903 -1084 937
rect 1084 903 1192 937
rect -1192 891 1192 903
rect -1192 841 -1134 891
rect -1192 -841 -1180 841
rect -1146 -841 -1134 841
rect 1134 841 1192 891
rect -1192 -891 -1134 -841
rect 1134 -841 1146 841
rect 1180 -841 1192 841
rect 1134 -891 1192 -841
rect -1192 -903 1192 -891
rect -1192 -937 -1084 -903
rect 1084 -937 1192 -903
rect -1192 -949 1192 -937
<< mvpsubdiffcont >>
rect -1084 903 1084 937
rect -1180 -841 -1146 841
rect 1146 -841 1180 841
rect -1084 -937 1084 -903
<< poly >>
rect -1000 799 1000 815
rect -1000 765 -984 799
rect 984 765 1000 799
rect -1000 727 1000 765
rect -1000 489 1000 527
rect -1000 455 -984 489
rect 984 455 1000 489
rect -1000 439 1000 455
rect -1000 381 1000 397
rect -1000 347 -984 381
rect 984 347 1000 381
rect -1000 309 1000 347
rect -1000 71 1000 109
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -109 1000 -71
rect -1000 -347 1000 -309
rect -1000 -381 -984 -347
rect 984 -381 1000 -347
rect -1000 -397 1000 -381
rect -1000 -455 1000 -439
rect -1000 -489 -984 -455
rect 984 -489 1000 -455
rect -1000 -527 1000 -489
rect -1000 -765 1000 -727
rect -1000 -799 -984 -765
rect 984 -799 1000 -765
rect -1000 -815 1000 -799
<< polycont >>
rect -984 765 984 799
rect -984 455 984 489
rect -984 347 984 381
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -381 984 -347
rect -984 -489 984 -455
rect -984 -799 984 -765
<< locali >>
rect -1180 903 -1084 937
rect 1084 903 1180 937
rect -1180 841 -1146 903
rect 1146 841 1180 903
rect -1000 765 -984 799
rect 984 765 1000 799
rect -1046 715 -1012 731
rect -1046 523 -1012 539
rect 1012 715 1046 731
rect 1012 523 1046 539
rect -1000 455 -984 489
rect 984 455 1000 489
rect -1000 347 -984 381
rect 984 347 1000 381
rect -1046 297 -1012 313
rect -1046 105 -1012 121
rect 1012 297 1046 313
rect 1012 105 1046 121
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -121 -1012 -105
rect -1046 -313 -1012 -297
rect 1012 -121 1046 -105
rect 1012 -313 1046 -297
rect -1000 -381 -984 -347
rect 984 -381 1000 -347
rect -1000 -489 -984 -455
rect 984 -489 1000 -455
rect -1046 -539 -1012 -523
rect -1046 -731 -1012 -715
rect 1012 -539 1046 -523
rect 1012 -731 1046 -715
rect -1000 -799 -984 -765
rect 984 -799 1000 -765
rect -1180 -903 -1146 -841
rect 1146 -903 1180 -841
rect -1180 -937 -1084 -903
rect 1084 -937 1180 -903
<< viali >>
rect -984 765 984 799
rect -1046 539 -1012 715
rect 1012 539 1046 715
rect -984 455 984 489
rect -984 347 984 381
rect -1046 121 -1012 297
rect 1012 121 1046 297
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -297 -1012 -121
rect 1012 -297 1046 -121
rect -984 -381 984 -347
rect -984 -489 984 -455
rect -1046 -715 -1012 -539
rect 1012 -715 1046 -539
rect -984 -799 984 -765
<< metal1 >>
rect -996 799 996 805
rect -996 765 -984 799
rect 984 765 996 799
rect -996 759 996 765
rect -1052 715 -1006 727
rect -1052 539 -1046 715
rect -1012 539 -1006 715
rect -1052 527 -1006 539
rect 1006 715 1052 727
rect 1006 539 1012 715
rect 1046 539 1052 715
rect 1006 527 1052 539
rect -996 489 996 495
rect -996 455 -984 489
rect 984 455 996 489
rect -996 449 996 455
rect -996 381 996 387
rect -996 347 -984 381
rect 984 347 996 381
rect -996 341 996 347
rect -1052 297 -1006 309
rect -1052 121 -1046 297
rect -1012 121 -1006 297
rect -1052 109 -1006 121
rect 1006 297 1052 309
rect 1006 121 1012 297
rect 1046 121 1052 297
rect 1006 109 1052 121
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -121 -1006 -109
rect -1052 -297 -1046 -121
rect -1012 -297 -1006 -121
rect -1052 -309 -1006 -297
rect 1006 -121 1052 -109
rect 1006 -297 1012 -121
rect 1046 -297 1052 -121
rect 1006 -309 1052 -297
rect -996 -347 996 -341
rect -996 -381 -984 -347
rect 984 -381 996 -347
rect -996 -387 996 -381
rect -996 -455 996 -449
rect -996 -489 -984 -455
rect 984 -489 996 -455
rect -996 -495 996 -489
rect -1052 -539 -1006 -527
rect -1052 -715 -1046 -539
rect -1012 -715 -1006 -539
rect -1052 -727 -1006 -715
rect 1006 -539 1052 -527
rect 1006 -715 1012 -539
rect 1046 -715 1052 -539
rect 1006 -727 1052 -715
rect -996 -765 996 -759
rect -996 -799 -984 -765
rect 984 -799 996 -765
rect -996 -805 996 -799
<< properties >>
string FIXED_BBOX -1163 -920 1163 920
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 10.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
