magic
tech sky130A
magscale 1 2
timestamp 1717253844
<< pwell >>
rect -201 -18582 201 18582
<< psubdiff >>
rect -165 18512 -69 18546
rect 69 18512 165 18546
rect -165 18450 -131 18512
rect 131 18450 165 18512
rect -165 -18512 -131 -18450
rect 131 -18512 165 -18450
rect -165 -18546 -69 -18512
rect 69 -18546 165 -18512
<< psubdiffcont >>
rect -69 18512 69 18546
rect -165 -18450 -131 18450
rect 131 -18450 165 18450
rect -69 -18546 69 -18512
<< xpolycontact >>
rect -35 17984 35 18416
rect -35 -18416 35 -17984
<< xpolyres >>
rect -35 -17984 35 17984
<< locali >>
rect -165 18512 -69 18546
rect 69 18512 165 18546
rect -165 18450 -131 18512
rect 131 18450 165 18512
rect -165 -18512 -131 -18450
rect 131 -18512 165 -18450
rect -165 -18546 -69 -18512
rect 69 -18546 165 -18512
<< viali >>
rect -19 18001 19 18398
rect -19 -18398 19 -18001
<< metal1 >>
rect -25 18398 25 18410
rect -25 18001 -19 18398
rect 19 18001 25 18398
rect -25 17989 25 18001
rect -25 -18001 25 -17989
rect -25 -18398 -19 -18001
rect 19 -18398 25 -18001
rect -25 -18410 25 -18398
<< properties >>
string FIXED_BBOX -148 -18529 148 18529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 180.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 1.029meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
